* NGSPICE file created from adc_array_matrix_flat.ext - technology: sky130A

.subckt adc_array_matrix_flat sample_n sample vcom row_n[0] row_n[1] row_n[2] row_n[3]
+ row_n[4] row_n[5] row_n[6] row_n[7] row_n[8] row_n[9] row_n[10] row_n[11] row_n[12]
+ row_n[13] row_n[14] row_n[15] row_n[16] row_n[17] row_n[18] row_n[19] row_n[20]
+ row_n[21] row_n[22] row_n[23] row_n[24] row_n[25] row_n[26] row_n[27] row_n[28]
+ row_n[29] row_n[30] row_n[31] en_n_bit[2] en_n_bit[1] en_n_bit[0] sw_n sw ctop analog_in
+ col_n[0] col_n[1] col_n[2] col_n[3] col_n[4] col_n[5] col_n[6] col_n[7] col_n[8]
+ col_n[9] col_n[10] col_n[11] col_n[12] col_n[13] col_n[14] col_n[15] colon_n[0]
+ colon_n[1] colon_n[2] colon_n[3] colon_n[4] colon_n[5] colon_n[6] colon_n[7] colon_n[8]
+ colon_n[9] colon_n[10] colon_n[11] colon_n[12] colon_n[13] colon_n[14] colon_n[15]
+ VSS VDD
X0 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=4.352e+14p ps=2.01194e+09u w=420000u l=150000u
X3 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=1.72952e+14p ps=1.48678e+09u w=800000u l=150000u
X4 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=7.7469e+13p pd=8.687e+08u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X6 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X7 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X8 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X9 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=1.4756e+14p ps=1.3209e+09u w=800000u l=150000u
X10 VSS col_n[0] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X11 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X12 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X13 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X14 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X15 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X16 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X17 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X18 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X19 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X20 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X21 VSS col_n[11] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X22 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X23 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X24 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X25 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X26 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X27 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X28 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X29 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X30 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X31 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X32 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X33 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X34 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X35 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X36 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X37 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X38 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X39 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X40 VSS col_n[8] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X41 VDD sample adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X42 VDD VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X43 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X44 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X45 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X46 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X47 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X48 VSS col_n[1] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X49 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X50 VSS col_n[13] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X51 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X52 VSS col_n[7] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X53 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X54 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X55 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X56 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X57 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X58 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X59 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X60 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X61 VSS col_n[14] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X62 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X63 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X64 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X65 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X66 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X67 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X68 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X69 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X70 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X71 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X72 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X73 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X74 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X75 VDD VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X76 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X77 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X78 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X79 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X80 VSS col_n[6] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X81 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X82 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X83 VSS col_n[2] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X84 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X85 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X86 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X87 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X88 VSS col_n[5] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X89 VSS sample_n adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X90 vcom VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X91 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X92 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X93 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X94 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X95 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X96 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X97 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X98 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X99 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X100 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X101 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X102 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X103 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X104 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X105 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X106 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X107 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X108 VSS col_n[12] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X109 VSS col_n[4] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X110 VSS col_n[0] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X111 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X112 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X113 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X114 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X115 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X116 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X117 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X118 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X119 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X120 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X121 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X122 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X123 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X124 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X125 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X126 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X127 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X128 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X129 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X130 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X131 vcom VSS adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X132 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X133 vcom VSS adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X134 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X135 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X136 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X137 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X138 VSS sample adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X139 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X140 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X141 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X142 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X143 VSS col_n[15] adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X144 VSS col_n[15] adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X145 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X146 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X147 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X148 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X149 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X150 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X151 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X153 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X154 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X155 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X156 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X157 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X158 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X159 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X160 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X161 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X162 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X163 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X164 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X165 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X166 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X167 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X168 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X169 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X170 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X171 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X172 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X173 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X174 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X175 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X176 VSS col_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X177 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X178 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X179 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X180 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X181 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X182 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X183 VSS VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X184 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X185 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X186 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X187 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X188 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X189 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X190 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X191 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X192 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X193 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X194 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X195 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X196 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X197 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X198 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X199 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X200 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X201 VSS col_n[11] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X202 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X203 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X204 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X205 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X206 VSS col_n[11] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X207 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X208 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X209 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X210 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X211 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X212 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X213 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X214 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X215 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X216 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X217 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X218 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X219 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X220 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X221 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X222 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X223 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X224 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X225 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X226 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X227 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X228 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X229 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X230 VSS VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X231 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X232 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X233 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X234 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X235 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X236 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X237 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X238 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X239 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X240 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X241 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X242 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X243 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X244 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X245 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X246 VSS col_n[1] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X247 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X248 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X249 VSS col_n[4] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X250 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X251 VSS col_n[7] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X252 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X253 VSS col_n[3] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X254 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X255 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X256 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X257 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X258 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X259 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X260 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X261 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X262 VDD colon_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X263 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X264 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X265 VSS col_n[9] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X266 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X267 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X268 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X269 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X270 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X271 VSS VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X272 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X273 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X274 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X275 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X276 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X277 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X278 VSS col_n[6] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X279 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X280 VDD VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X281 VSS col_n[2] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X282 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X283 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X284 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X285 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X286 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X287 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X288 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X289 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X290 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X291 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X292 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X293 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X294 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X295 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X296 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X297 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X298 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X299 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X300 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X301 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X302 VSS sample_n adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X303 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X304 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X305 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X306 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X307 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X308 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X309 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X310 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X311 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X312 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X313 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X314 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X315 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X316 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X317 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X318 VSS col_n[11] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X319 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X320 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X321 VSS col_n[10] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X322 VSS col_n[10] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X323 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X324 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X325 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X326 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X327 VSS col_n[4] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X328 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X329 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X330 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X331 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X332 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X333 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X334 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X335 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X336 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X337 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X338 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X339 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X340 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X341 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X342 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X343 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X344 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X345 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X346 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X347 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X348 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X349 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X350 VSS col_n[8] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X351 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X352 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X353 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X354 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X355 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X356 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X357 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X358 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X359 vcom VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X360 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X361 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X362 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X363 vcom VSS adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X364 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X365 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X366 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X367 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X368 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X369 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X370 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X371 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X372 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X373 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X374 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X375 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X376 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X377 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X378 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X379 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X380 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X381 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X382 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X383 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X384 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X385 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X386 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X387 vcom VSS adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X388 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X389 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X390 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X391 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X392 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X393 VDD sample adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X394 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X395 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X396 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X397 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X398 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X399 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X400 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X401 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X402 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X403 VSS col_n[5] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X404 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X405 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X406 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X407 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X408 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X409 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X410 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X411 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X412 VSS col_n[12] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X413 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X414 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X415 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X416 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X417 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X418 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X419 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X420 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X421 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X422 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X423 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X424 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X425 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X426 VSS col_n[1] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X427 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X428 VSS col_n[4] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X429 VSS col_n[0] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X430 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X431 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X432 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X433 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X434 VSS sample_n adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X435 VSS col_n[3] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X436 VSS col_n[7] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X437 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X438 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X439 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X440 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X441 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X442 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X443 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X444 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X445 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X446 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X447 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X448 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X449 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X450 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X451 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X452 VSS VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X453 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X454 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X455 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X456 VSS VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X457 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X458 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X459 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X460 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X461 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X462 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X463 VSS col_n[2] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X464 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X465 VSS col_n[6] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X466 VDD VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X467 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X468 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X469 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X470 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X471 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X472 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X473 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X474 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X475 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X476 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X477 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X478 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X479 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X480 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X481 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X482 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X483 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X484 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X485 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X486 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X487 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X488 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X489 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X490 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X491 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X492 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X493 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X494 VSS col_n[13] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X495 VSS col_n[13] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X496 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X497 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X498 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X499 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X500 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X501 VSS col_n[6] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X502 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X503 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X504 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X505 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X506 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X507 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X508 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X509 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X510 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X511 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X512 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X513 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X514 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X515 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X516 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X517 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X518 VSS col_n[11] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X519 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X520 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X521 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X522 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X523 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X524 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X525 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X526 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X527 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X528 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X529 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X530 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X531 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X532 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X533 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X534 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X535 VSS col_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X536 VSS VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X537 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X538 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X539 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X540 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X541 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X542 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X543 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X544 VSS col_n[14] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X545 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X546 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X547 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X548 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X549 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X550 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X551 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X552 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X553 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X554 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X555 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X556 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X557 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X558 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X559 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X560 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X561 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X562 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X563 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X564 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X565 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X566 VDD VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X567 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X568 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X569 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X570 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X571 VSS col_n[1] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X572 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X573 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X574 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X575 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X576 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X577 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X578 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X579 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X580 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X581 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X582 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X583 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X584 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X585 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X586 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X587 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X588 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X589 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X590 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X591 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X592 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X593 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X594 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X595 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X596 VSS col_n[11] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X597 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X598 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X599 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X600 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X601 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X602 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X603 VSS col_n[2] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X604 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X605 VSS col_n[5] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X606 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X607 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X608 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X609 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X610 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X611 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X612 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X613 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X614 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X615 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X616 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X617 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X618 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X619 VSS col_n[14] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X620 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X621 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X622 VSS col_n[1] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X623 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X624 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X625 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X626 VSS col_n[4] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X627 VSS col_n[0] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X628 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X629 VDD VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X630 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X631 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X632 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X633 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X634 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X635 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X636 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X637 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X638 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X639 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X640 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X641 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X642 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X643 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X644 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X645 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X646 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X647 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X648 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X649 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X650 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X651 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X652 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X653 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X654 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X655 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X656 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X657 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X658 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X660 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X661 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X662 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X663 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X664 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X665 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X666 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X667 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X668 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X669 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X670 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X671 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X672 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X673 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X674 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X675 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X676 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X677 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X678 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X679 vcom VSS adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X680 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X681 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X682 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X683 VSS col_n[6] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X684 vcom VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X685 VSS col_n[2] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X686 vcom VSS adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X687 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X688 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X689 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X690 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X691 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X692 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X693 VSS col_n[15] adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X694 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X695 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X696 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X697 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X698 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X699 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X700 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X701 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X702 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X703 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X704 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X705 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X706 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X707 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X708 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X709 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X710 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X711 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X712 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X713 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X714 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X715 VSS VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X716 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X717 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X718 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X719 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X720 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X721 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X722 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X723 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X724 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X725 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X726 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X727 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X728 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X729 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X730 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X731 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X732 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X733 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X734 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X735 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X736 VSS col_n[9] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X737 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X738 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X739 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X740 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X741 VDD sample_n adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X742 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X743 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X744 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X745 VSS VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X746 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X747 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X748 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X749 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X750 vcom VSS adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X751 VSS col_n[15] adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X752 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X753 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X754 VSS col_n[1] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X755 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X756 VSS col_n[11] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X757 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X758 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X759 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X760 VSS col_n[11] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X761 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X762 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X763 VSS col_n[3] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X764 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X765 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X766 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X767 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X768 VSS col_n[7] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X769 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X770 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X771 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X772 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X773 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X774 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X775 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X776 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X777 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X778 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X779 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X780 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X781 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X782 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X783 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X784 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X785 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X786 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X787 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X788 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X789 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X790 VSS col_n[2] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X791 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X792 VSS col_n[6] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X793 VSS sample_n adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X794 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X795 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X796 VSS col_n[5] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X797 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X798 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X799 VSS col_n[14] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X800 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X801 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X802 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X803 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X804 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X805 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X806 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X807 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X808 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X809 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X810 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X811 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X812 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X813 VSS col_n[0] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X814 VDD VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X815 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X816 VSS col_n[9] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X817 VSS col_n[4] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X818 VSS VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X819 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X820 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X821 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X822 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X823 VSS col_n[11] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X824 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X825 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X826 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X827 VSS col_n[6] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X828 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X829 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X830 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X831 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X832 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X833 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X834 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X835 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X836 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X837 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X838 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X839 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X840 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X841 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X842 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X843 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X844 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X845 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X846 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X847 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X848 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X849 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X850 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X851 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X852 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X853 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X854 VSS col_n[4] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X855 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X856 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X857 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X858 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X859 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X860 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X861 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X862 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X863 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X864 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X865 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X866 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X867 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X868 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X869 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X870 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X871 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X872 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X873 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X874 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X875 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X876 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X877 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X878 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X879 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X880 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X881 VSS col_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X882 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X883 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X884 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X885 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X886 VSS col_n[6] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X887 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X888 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X889 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X890 VDD sample_n adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X891 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X892 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X893 VSS col_n[12] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X894 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X895 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X896 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X897 VSS col_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X898 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X899 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X900 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X901 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X902 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X903 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X904 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X905 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X906 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X907 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X908 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X909 VSS col_n[10] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X910 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X911 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X912 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X913 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X914 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X915 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X916 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X917 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X918 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X919 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X920 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X921 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X922 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X923 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X924 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X925 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X926 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X927 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X928 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X929 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X930 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X931 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X932 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X933 VSS col_n[15] adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X934 VSS col_n[15] adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X935 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X936 ctop sw_n analog_in VDD sky130_fd_pr__pfet_01v8 ad=5.9e+11p pd=3.18e+06u as=5.8e+11p ps=5.16e+06u w=1e+06u l=1e+06u
X937 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X938 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X939 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X940 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X941 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X942 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X943 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X944 VDD sample adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X945 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X946 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X947 vcom VSS adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X948 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X949 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X950 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X951 VSS col_n[1] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X952 VSS col_n[10] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X953 VSS col_n[0] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X954 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X955 VSS col_n[7] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X956 VSS col_n[3] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X957 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X958 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X959 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X960 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X961 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X962 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X963 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X964 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X965 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X966 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X967 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X968 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X969 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X970 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X971 VSS col_n[12] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X972 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X973 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X974 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X975 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X976 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X977 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X978 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X979 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X980 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X981 VSS col_n[2] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X982 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X983 vcom VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X984 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X985 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X986 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X987 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X988 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X989 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X990 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X991 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X992 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X993 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X994 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X995 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X996 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X997 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X998 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X999 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1000 VSS col_n[9] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1001 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X1002 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1003 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1004 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1005 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1006 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1007 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1008 VSS col_n[6] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1009 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1010 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1011 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1012 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1013 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1014 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1015 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1016 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1017 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1018 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1019 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1020 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1021 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1022 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1023 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1024 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1025 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1026 VSS col_n[7] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1027 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1028 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1029 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1030 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1031 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1032 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1033 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1034 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1035 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1036 VSS col_n[4] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1037 VSS col_n[0] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1038 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1039 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1040 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1041 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1042 VDD VSS adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1043 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1044 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1045 VSS col_n[13] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1046 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1047 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1048 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1049 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1050 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1051 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1052 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1053 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1054 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1055 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1056 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1057 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1058 VSS VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1059 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1060 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1061 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1062 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1063 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1064 VSS col_n[8] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1065 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1066 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1067 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1068 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1069 vcom VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1070 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1071 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1072 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1073 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1074 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1075 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1076 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1077 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1078 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1079 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1080 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1081 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1082 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1083 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1084 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1085 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1086 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1087 VDD sample adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1088 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1089 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1090 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1091 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1092 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1093 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1094 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1095 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1096 VSS col_n[14] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1097 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1098 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1099 VSS col_n[13] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1100 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1101 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1102 vcom VSS adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1103 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1104 VDD VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1105 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1106 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1107 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1108 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1109 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1110 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1111 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1112 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1113 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1114 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1115 VSS col_n[5] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1116 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1117 VSS col_n[10] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1118 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1119 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1120 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1121 VSS col_n[10] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1122 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1123 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1124 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1125 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1126 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1127 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1128 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1129 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1130 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1131 VSS col_n[0] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1132 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1133 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1134 VSS col_n[4] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1135 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1136 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1137 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1138 VSS col_n[3] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1139 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1140 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1141 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1142 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1143 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1144 VSS col_n[12] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1145 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1146 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1147 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1148 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1149 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1150 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1151 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1152 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1153 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1154 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1155 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1156 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1157 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1158 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1159 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1160 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1161 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1162 VDD VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1163 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1164 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1165 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1166 VDD VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1167 VSS col_n[2] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1168 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1169 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1170 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1171 VSS col_n[4] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1172 VSS col_n[15] adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1173 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1174 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1175 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1176 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1177 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1178 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1179 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1180 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1181 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1182 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1183 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1184 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1185 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1186 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1187 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1188 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1189 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1190 VDD VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1191 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1192 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1193 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1194 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1195 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1196 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1197 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1198 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1199 VSS col_n[6] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1200 VSS col_n[2] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1201 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1202 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1203 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1204 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1205 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1206 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1207 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1208 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1209 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1210 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1211 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1212 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1213 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1214 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1215 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1216 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1217 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1218 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1219 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1220 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1221 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1222 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1223 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1224 VSS col_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1225 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1226 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1227 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1228 VSS col_n[4] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1229 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1230 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1231 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1232 VDD sample_n adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1233 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1234 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1235 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1236 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1237 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1238 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1239 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1240 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1241 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1242 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1243 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1244 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1245 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1246 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1247 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1248 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1249 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1250 vcom VSS adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1251 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1252 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1253 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1254 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1255 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1256 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1257 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1258 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1259 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1260 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1261 VSS col_n[1] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1262 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1263 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1264 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1265 VSS col_n[13] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1266 VSS col_n[13] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1267 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1268 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1269 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1270 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1271 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1272 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1273 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1274 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1275 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1276 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1277 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1278 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1279 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1280 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1281 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1282 VDD sample adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1283 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1284 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1285 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1286 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1287 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1288 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1289 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1290 VSS col_n[9] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1291 vcom VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1292 VSS VSS adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1293 VSS col_n[5] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1294 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1295 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1296 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1297 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1298 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1299 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1300 VSS VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1301 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1302 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1303 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1304 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1305 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1306 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1307 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1308 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1309 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1310 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1311 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1312 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1313 VSS col_n[0] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1314 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1315 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1316 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1317 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1318 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1319 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1320 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1321 VSS col_n[6] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1322 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1323 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1324 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1325 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1326 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1327 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1328 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1329 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1330 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1331 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1332 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1333 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1334 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1335 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1336 vcom VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1337 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1338 VSS col_n[4] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1339 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1340 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1341 VSS col_n[7] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1342 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1343 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1344 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1345 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1346 VSS col_n[10] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1347 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1348 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1349 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1350 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1351 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1352 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1353 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1354 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1355 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1356 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1357 VSS col_n[11] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1358 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1359 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1360 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1361 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1362 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1363 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1364 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1365 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1366 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1367 VSS col_n[5] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1368 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1369 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1370 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1371 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1372 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1373 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1374 VSS col_n[2] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1375 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1376 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1377 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1378 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1379 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1380 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1381 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1382 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1383 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1384 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1385 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1386 VDD VSS adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1387 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1388 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1389 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1390 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1391 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1392 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1393 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1394 VSS col_n[14] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1395 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1396 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1397 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1398 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1399 VSS VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1400 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1401 VSS VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1402 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1403 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1404 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1405 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1406 VDD VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1407 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1408 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1409 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1410 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1411 VSS sample adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1412 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1413 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1414 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1415 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1416 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1417 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1418 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1419 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1420 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1421 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1422 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1423 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1424 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1425 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1426 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1427 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1428 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1429 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1430 VSS col_n[12] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1431 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1432 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1433 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1434 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1435 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1436 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1437 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1438 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1439 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1440 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1441 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1442 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1443 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1444 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1445 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1446 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1447 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1448 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1449 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1450 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1451 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1452 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1453 VSS col_n[3] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1454 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1455 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1456 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1457 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1458 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1459 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1460 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1461 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1462 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1463 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1464 VSS VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1465 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1466 VSS VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1467 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1468 VSS col_n[15] adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1469 VSS col_n[15] adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1470 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1471 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1472 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1473 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1474 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1475 VSS col_n[2] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1476 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1477 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1478 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1479 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1480 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1481 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1482 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1483 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1484 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1485 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1486 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1487 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1488 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1489 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1490 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1491 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1492 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1493 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1494 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1495 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1496 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1497 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1498 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1499 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1500 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1501 VSS col_n[0] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1502 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1503 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1504 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1505 VSS col_n[6] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 VSS col_n[2] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1507 VSS col_n[13] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1508 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1509 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1510 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1511 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1512 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1513 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1514 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1515 VSS col_n[8] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1516 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1517 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1518 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1519 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1520 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1521 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1522 VDD colon_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1523 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1524 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1525 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1526 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1527 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1528 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1529 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1530 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1531 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1532 VDD colon_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1533 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1534 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1535 VSS col_n[11] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1536 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1537 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1538 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1539 VSS col_n[4] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1540 VSS col_n[0] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1541 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1542 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1543 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1544 VSS col_n[7] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1545 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1546 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1547 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1548 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1549 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1550 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1551 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1552 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1553 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1554 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1555 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1556 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1557 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1558 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1559 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1560 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1561 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1562 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1563 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1564 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1565 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1566 vcom VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1567 vcom VSS adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1568 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1569 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1570 VSS col_n[2] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1571 VDD sample_n adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1572 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1573 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1574 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1575 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1576 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1577 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1578 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1579 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1580 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1581 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1582 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1583 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1584 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1585 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1586 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1587 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1588 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1589 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1590 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1591 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1592 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1593 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1594 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1595 VSS col_n[9] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1596 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1597 VSS VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1598 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1599 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1600 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1601 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1602 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1603 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1604 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1605 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1606 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1607 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1608 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1609 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1610 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1611 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1612 VDD VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1613 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1614 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1615 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1616 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1617 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1618 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1619 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1620 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1621 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1622 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1623 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1624 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1625 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1626 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1627 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1628 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1629 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1630 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1631 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1632 VSS col_n[3] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1633 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1634 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1635 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1636 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1637 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1638 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1639 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1640 VSS col_n[14] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1641 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1642 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1643 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1644 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1645 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1646 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1647 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1648 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1649 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1650 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1651 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1652 VDD VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1653 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1654 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1655 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1656 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1657 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1658 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1659 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1660 VSS col_n[10] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1661 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1662 VSS col_n[10] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1663 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1664 VSS col_n[4] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1665 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1666 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1667 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1668 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1669 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1670 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1671 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1672 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1673 VDD colon_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1674 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1675 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1676 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1677 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1678 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1679 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1680 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1681 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1682 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1683 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1684 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1685 VSS col_n[6] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1686 VSS col_n[2] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1687 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1688 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1689 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1690 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1691 VSS col_n[5] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1692 VSS col_n[8] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1693 VSS sample_n adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1694 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1695 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1696 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1697 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1698 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1699 vcom VSS adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1700 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1701 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1702 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1703 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1704 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1705 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1706 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1707 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1708 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1709 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1710 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1711 VSS col_n[15] adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1712 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1713 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1714 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1715 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1716 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1717 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1718 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1719 VSS col_n[7] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1720 VSS col_n[3] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1721 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1722 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1723 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1724 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1725 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1726 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1727 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1728 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1729 VSS col_n[0] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1730 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X1731 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1732 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1733 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1734 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1735 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1736 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1737 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1738 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1739 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1740 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1741 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1742 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1743 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1744 VSS col_n[12] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1746 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1747 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint2 en_n_bit[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1748 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1749 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1750 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1751 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1752 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1753 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1754 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1755 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1756 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1757 VSS sample adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1758 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1759 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1760 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1761 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1762 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1763 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1764 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1765 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1766 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1767 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1768 VSS VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1769 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1770 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1771 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1772 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1773 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1774 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1775 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1776 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1777 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1778 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1779 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1780 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1781 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1782 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1783 vcom VSS adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1784 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1785 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1786 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1787 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1788 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1789 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1790 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1791 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1792 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1793 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1794 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1795 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1796 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1797 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1798 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1799 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1800 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1801 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1802 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1803 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1804 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1805 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1806 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1807 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1808 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1809 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1810 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1811 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1812 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1813 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1814 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1815 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1816 VSS col_n[14] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1817 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1818 VSS col_n[14] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1819 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1820 VSS col_n[13] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 VSS col_n[13] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1822 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1823 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1824 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1825 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1826 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1827 VSS col_n[6] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1828 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1829 VSS col_n[0] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1830 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1831 VDD VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1832 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1833 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1834 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1835 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1836 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1837 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1838 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1839 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1840 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1841 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1842 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1843 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1844 VSS col_n[9] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1845 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1846 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1847 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1848 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1849 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1850 VSS col_n[11] adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1851 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1852 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1853 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1854 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1855 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1856 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1857 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1858 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1859 VSS VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1860 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1861 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1862 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1863 VSS col_n[4] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1864 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1865 VSS col_n[0] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1866 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1867 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1868 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1869 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1870 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1871 VSS col_n[7] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1872 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1873 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1874 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1875 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1876 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1877 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1878 VDD colon_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1879 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1880 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1881 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1882 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1883 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1884 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1885 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1886 VDD colon_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1887 VSS col_n[2] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1888 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1889 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1890 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1891 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1892 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1893 VSS col_n[6] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1894 VSS col_n[5] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1895 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1896 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1897 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1898 vcom VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1899 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1900 VSS VSS adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1901 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1902 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1903 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1904 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1905 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1906 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1907 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1908 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1909 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1910 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X1911 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1912 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X1913 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1914 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1915 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1916 VSS col_n[10] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1917 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1918 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1919 VSS sample_n adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1920 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1921 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1922 VSS col_n[0] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1923 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1924 VDD sample_n adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1925 VSS col_n[11] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1926 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1927 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1928 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1929 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1930 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1931 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1932 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1933 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1934 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1935 VDD VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1936 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1937 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1938 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1939 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1940 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1941 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1942 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1943 VSS col_n[14] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1944 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1945 VSS col_n[1] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1946 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1947 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1948 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1949 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1950 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1951 VSS col_n[7] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1952 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1953 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1954 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1955 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1956 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1957 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X1958 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1959 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1960 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1961 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1962 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1963 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1964 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1965 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1966 VDD VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1967 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1968 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1969 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1970 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1971 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1972 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1973 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1974 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1975 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1976 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1977 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1978 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1979 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1980 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1981 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1982 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X1983 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1984 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1985 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1986 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1987 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1988 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1989 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X1990 VDD VSS adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1991 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X1992 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1993 VSS col_n[12] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X1994 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X1995 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1996 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X1997 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X1998 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X1999 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2000 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2001 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2002 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2003 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2004 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2005 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2006 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2007 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2008 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2009 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2010 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2011 VSS col_n[9] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2012 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2013 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X2014 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2015 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2016 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2017 VSS col_n[9] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2018 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2019 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2020 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2021 VSS col_n[6] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2022 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2023 VSS col_n[2] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2024 VSS VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2025 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2026 VSS VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2027 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2028 VSS col_n[8] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2029 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2030 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2031 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2032 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2033 VSS col_n[15] adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2034 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2035 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2036 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2037 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2038 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2039 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2040 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2041 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2042 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2043 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2044 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2045 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2046 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2047 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2048 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2049 VSS col_n[4] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2050 VSS col_n[0] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2051 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2052 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2053 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2054 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2055 VSS col_n[7] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2056 VSS sample_n adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2057 VSS col_n[3] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2058 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2059 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2060 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2061 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2062 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2063 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2064 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2065 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2066 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2067 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2068 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2069 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2070 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2071 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2072 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2073 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2074 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2075 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2076 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2077 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2078 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2079 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2080 VSS col_n[13] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2081 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2082 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2083 VSS col_n[5] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2084 vcom VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2085 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2086 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2087 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2088 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2089 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2090 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2091 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2092 VSS VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2093 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2094 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2095 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2096 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2097 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2098 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2099 VSS col_n[11] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2100 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2101 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2102 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2103 VSS col_n[11] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2104 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2105 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2106 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2107 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2108 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2109 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2110 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2111 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2112 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2113 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2114 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2115 VSS sample adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2116 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2117 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2118 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2119 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2120 VSS sample_n adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2121 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2122 VSS VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2123 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2124 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2125 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2126 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2127 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2128 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2129 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2130 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2131 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2132 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2133 VSS col_n[14] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2134 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2135 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2136 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2137 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2138 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2139 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2140 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2141 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2142 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2143 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2144 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2145 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2146 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2147 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2148 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2149 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2150 VDD VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2151 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2152 VSS col_n[9] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2153 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2154 VSS col_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2155 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2156 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2157 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2158 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2159 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2160 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2161 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2162 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2163 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2164 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2165 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2166 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2167 VSS VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2168 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2169 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2170 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2171 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2172 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2173 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2174 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2175 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2176 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2177 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2178 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2179 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2180 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2181 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2182 VSS col_n[12] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2183 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2184 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2185 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2186 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2187 VSS col_n[12] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2188 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2189 vcom VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2190 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2191 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2192 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2193 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2194 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2195 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2196 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2197 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2198 VSS col_n[4] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2199 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2200 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2201 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2202 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2203 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2204 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2205 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2206 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2207 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2208 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2209 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2210 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2211 VSS VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2212 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2213 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2214 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2215 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2216 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2217 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2218 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2219 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2220 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2221 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2222 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2223 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2224 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2225 VSS col_n[14] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2226 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2227 VSS col_n[2] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2228 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2229 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2231 VSS col_n[6] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2232 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2233 VSS col_n[5] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2234 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2235 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2236 VSS col_n[8] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2237 VDD VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2238 VDD VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2239 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2240 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2241 VSS col_n[11] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2242 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2243 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2244 VDD colon_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2245 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2246 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2247 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2248 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2249 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2250 VSS col_n[10] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2251 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2252 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2253 VDD colon_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2254 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2255 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2256 VSS col_n[0] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2257 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2258 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2259 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2260 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2261 VSS col_n[4] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2262 VSS col_n[3] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2263 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2264 VSS col_n[7] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2265 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2266 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2267 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2268 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2269 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2270 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2271 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2272 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2273 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2274 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2275 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2276 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2277 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2278 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2279 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2280 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2281 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2282 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2283 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2284 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2285 VSS sample_n adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2287 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2288 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2289 vcom VSS adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2290 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2291 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2292 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2293 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2294 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2295 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2296 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2297 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2298 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2299 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2300 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2301 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2302 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2303 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2304 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2305 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2306 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2307 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2308 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2309 VDD VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2310 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2311 VSS col_n[12] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2312 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2313 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2314 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2315 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2316 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2317 VSS col_n[5] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2318 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2319 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2320 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2321 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2322 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2323 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2324 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2325 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2326 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2327 VDD VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2328 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2329 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2330 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2331 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2332 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2333 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2334 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2335 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2336 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2337 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2338 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2339 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2340 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2341 VSS col_n[9] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2342 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2343 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2344 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2345 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2346 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2347 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2348 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2349 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2350 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2351 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2352 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2353 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2354 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2355 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X2356 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2357 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2358 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2359 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2360 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2361 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2362 analog_in sw_n ctop VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2363 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2364 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2365 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2366 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2367 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2368 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2369 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2370 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2371 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2372 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2373 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2374 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2375 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2376 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2377 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2378 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2379 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2380 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2381 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2382 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2383 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2384 VSS col_n[4] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2385 VSS col_n[0] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2386 VSS col_n[14] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2387 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2388 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2389 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2390 VSS col_n[14] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2391 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2392 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2393 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2394 VSS col_n[13] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2395 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2396 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2397 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2398 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2399 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2400 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2401 VDD VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2402 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2403 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2404 VDD VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2405 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2406 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2407 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2408 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2409 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2410 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2411 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2412 VSS col_n[2] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2413 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2414 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2415 VSS col_n[5] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2416 VSS sample_n adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2417 VSS col_n[9] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2418 VSS col_n[8] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2419 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2420 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2421 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2422 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2423 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2424 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2425 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2426 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2427 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2428 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2429 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2430 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2431 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2432 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2433 vcom VSS adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2434 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2435 VSS col_n[1] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2436 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2437 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2438 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2439 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2440 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2441 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2442 VSS col_n[7] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2443 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2444 VSS col_n[3] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2445 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2446 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2447 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2448 VSS col_n[14] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2449 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2450 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2451 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2452 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2453 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2454 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2455 VDD VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2456 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2457 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2458 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2459 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2460 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2461 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2462 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2463 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2464 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2465 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2466 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2467 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2468 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2469 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2470 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2471 VSS sample adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2472 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2473 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2474 VSS col_n[7] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2475 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X2476 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2477 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2478 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2479 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2480 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2481 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2482 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2483 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2484 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2485 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2486 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2487 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2488 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2489 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2490 VSS VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2491 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2492 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2493 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2494 VSS col_n[12] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2495 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2496 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2497 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2498 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2499 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2500 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2501 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2502 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2503 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2504 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2505 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2506 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2507 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2508 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2509 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2510 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2511 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2512 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2513 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2514 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2515 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2516 VSS col_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2517 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2518 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2519 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2520 VSS VSS adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2521 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2522 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2523 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2524 VSS col_n[15] adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2525 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2526 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2527 VSS col_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2528 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2529 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2530 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2531 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2532 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2533 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2534 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2535 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2536 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2537 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2538 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2539 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2540 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2541 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2542 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2543 VDD VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2544 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2545 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2546 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2547 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2548 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2549 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2550 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2551 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2552 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2553 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2554 VSS col_n[6] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2555 VSS col_n[2] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2556 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2557 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2558 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2559 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2560 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2561 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2562 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2563 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2564 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2565 VDD VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2566 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2567 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2568 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2569 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2570 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2571 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2572 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2573 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2574 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2575 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2576 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2577 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2578 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2579 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2580 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2581 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2582 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2583 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2584 VSS col_n[12] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2585 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2586 VSS col_n[0] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2587 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2588 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2589 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2590 VSS col_n[4] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2591 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2592 VDD sample adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2593 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2594 VSS col_n[3] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2595 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X2596 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2597 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2598 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2599 VSS col_n[9] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2600 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2601 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2602 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2603 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2604 VSS col_n[9] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2605 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2606 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2607 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2608 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2609 VSS col_n[15] adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2610 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2611 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2612 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2613 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2614 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2615 vcom VSS adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2616 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2617 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2618 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2619 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2620 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2621 VSS col_n[2] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2622 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2623 VSS col_n[5] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2624 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2625 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2626 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2627 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2628 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2629 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2630 VDD VSS adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2631 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2632 VSS col_n[1] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2633 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2634 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2635 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2636 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2637 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2638 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2639 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2640 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2641 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2642 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2643 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2644 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2645 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2646 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2647 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2648 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2649 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2650 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2651 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2652 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2653 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2654 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2655 VSS col_n[9] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2656 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2657 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2658 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2659 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2660 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2661 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2662 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2663 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2664 VSS VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2665 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2666 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2667 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2668 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2669 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2670 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2671 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2672 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2673 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2674 VSS col_n[11] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2675 VSS col_n[11] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2676 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2677 VSS col_n[3] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2678 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2679 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2680 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2681 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2682 VSS col_n[7] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2683 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2684 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2685 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2686 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2687 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2688 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2689 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2690 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2691 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2692 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2693 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2694 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2695 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2696 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2697 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2698 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2699 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2700 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2701 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2702 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2703 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2704 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2705 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2706 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2707 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2708 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2709 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2710 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2711 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2712 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2713 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2714 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2715 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2716 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2717 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2718 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2719 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2720 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2721 VSS sample adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2722 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2723 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2724 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2725 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2726 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2727 VSS col_n[10] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2728 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2729 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2730 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2731 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2732 VSS col_n[9] adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2733 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2734 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2735 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2736 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2737 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2738 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2739 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2740 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2741 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X2742 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2743 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2744 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2745 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2746 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2747 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2748 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2749 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2750 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2751 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2752 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2753 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2754 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2755 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2756 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2757 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2758 VSS col_n[2] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2759 VSS col_n[12] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2760 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2761 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2762 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2763 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2764 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2765 VSS col_n[12] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2766 VSS col_n[8] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2767 VDD VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2768 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2769 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2770 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2771 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2772 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2773 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2774 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2775 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2776 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2777 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2778 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2779 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2780 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2781 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2782 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2783 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2784 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2785 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2786 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2787 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2788 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint1 en_n_bit[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2789 VSS col_n[0] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2790 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2791 VSS col_n[7] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2792 VSS col_n[3] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2793 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2794 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2795 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2796 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2797 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2798 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2799 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2800 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2801 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2802 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2803 VSS col_n[15] adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2804 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2805 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2806 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2807 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2808 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2809 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2810 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2811 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2812 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2813 vcom VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2814 VSS col_n[10] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2815 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2816 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2817 VSS col_n[5] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2818 vcom VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2819 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2820 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2821 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2822 VSS col_n[12] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2823 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2824 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2825 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2826 VSS col_n[7] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2827 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2828 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2829 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2830 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2831 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2832 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2833 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2834 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2835 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2836 adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2837 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2838 VSS VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2839 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2840 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2841 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2842 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2843 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2844 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2845 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2846 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2847 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2848 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2849 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2850 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2851 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2852 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2853 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2854 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2855 VSS VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2856 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X2857 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2858 VSS col_n[5] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2859 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2860 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2861 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2862 VSS VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2863 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2864 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2865 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2866 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2867 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2868 VDD en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2869 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2870 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2871 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2872 vcom VSS adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2873 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2874 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2875 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2876 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2877 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2878 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2879 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2880 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2881 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2882 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2883 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2884 VSS col_n[7] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2885 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint1 en_n_bit[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2886 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2887 VSS col_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2888 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2889 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2890 VDD sample_n adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2891 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2892 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2893 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2894 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2895 VSS col_n[13] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2896 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2897 VSS VSS adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2898 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2899 VSS col_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2900 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2901 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2902 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2903 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2904 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2905 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2906 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2907 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2908 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2909 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2910 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2911 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2912 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2913 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2914 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2915 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2916 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2917 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2918 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2919 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2920 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2921 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2922 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2923 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2924 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2925 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2926 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2927 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2928 VSS col_n[4] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2929 VSS col_n[0] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2930 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2931 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2932 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2933 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2934 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2935 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2936 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2937 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2938 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2939 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2940 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2941 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2942 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2943 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2944 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2945 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2946 VDD VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2947 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2948 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2949 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2950 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2951 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2952 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2953 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2954 VDD sample_n adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2955 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2956 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2957 VDD sample adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2958 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2959 VSS col_n[2] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2960 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2961 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X2962 VSS col_n[8] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2963 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X2964 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2965 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2966 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2967 VDD en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2968 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2969 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2970 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2971 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2972 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2973 VSS col_n[1] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2974 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2975 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2976 VSS col_n[13] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2977 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2978 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2979 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2980 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2981 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2982 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2983 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2984 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2985 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2986 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2987 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2988 VSS col_n[0] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X2989 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2990 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2991 VSS col_n[3] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2992 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X2993 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X2994 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2995 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X2996 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X2997 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2998 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X2999 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3000 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3001 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3002 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3003 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3004 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3005 vcom VSS adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3006 VSS col_n[10] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3007 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3008 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3009 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3010 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3011 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3012 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3013 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3014 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3015 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3016 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3017 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3018 VSS col_n[7] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3019 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3020 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3021 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3022 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3023 VSS VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3024 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X3025 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3026 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3027 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3028 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3029 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3030 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3031 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3032 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3033 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3034 VSS col_n[14] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3035 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3036 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3037 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3038 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3039 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3040 vcom VSS adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3041 VSS col_n[8] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3042 VDD VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3043 vcom VSS adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3044 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3045 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3046 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3047 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3048 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3049 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3050 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3051 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3052 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3053 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3054 VSS col_n[5] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3055 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3056 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3057 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3058 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3059 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3060 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3061 vcom VSS adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3062 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3063 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3064 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3065 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3066 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3067 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3068 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3069 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3070 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3071 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3072 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3073 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3074 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3075 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3076 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3077 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3078 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3079 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3080 adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3081 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3082 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3083 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3084 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3085 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3086 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3087 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3088 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3089 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3090 VSS sample adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3091 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3092 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3093 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3094 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3095 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3096 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3097 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3098 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3099 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3100 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3101 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3102 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3103 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3104 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3105 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3106 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3107 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3108 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3109 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3110 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3111 VSS col_n[15] adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3112 VDD sample_n adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3113 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3114 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3115 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3116 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3117 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3118 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3119 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3120 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3121 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3122 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3123 VSS col_n[0] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3124 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3125 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3126 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3127 VSS en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X3128 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3129 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3130 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3131 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3132 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3133 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3134 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3135 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3136 VDD VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3137 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3138 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3139 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3140 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3141 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3142 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3143 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3144 adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3145 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3146 VSS col_n[5] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3147 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3148 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3149 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3150 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3151 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3152 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3153 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3154 VSS col_n[13] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3155 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3156 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3157 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3158 VSS col_n[1] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3159 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3160 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3161 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3162 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3163 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3164 VSS VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3165 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3166 VSS col_n[3] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3167 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3168 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3169 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3170 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3171 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3172 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3173 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3174 vcom VSS adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3175 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3176 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3177 VSS col_n[5] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3178 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3179 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3180 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3181 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3182 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3183 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3184 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3185 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3186 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3187 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3188 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3189 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3190 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3191 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3192 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3193 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3194 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3195 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3196 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3197 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3198 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint2 en_n_bit[0] adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3199 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3200 VSS col_n[14] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3201 VSS col_n[7] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3202 VSS col_n[3] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3203 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3204 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3205 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3206 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3207 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3208 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3209 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3210 VSS en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3211 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3212 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3213 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3214 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3215 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3216 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3217 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3218 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3219 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3220 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3221 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3222 VSS col_n[9] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3223 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3224 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3225 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3226 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3227 VSS col_n[5] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3228 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3229 VDD sample_n adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3230 VSS VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3231 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3232 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3233 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3234 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3235 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3236 adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3237 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3238 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3239 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3240 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3241 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3242 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3243 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3244 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3245 VSS col_n[11] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3246 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3247 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3248 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3249 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3250 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3251 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3252 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3253 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3254 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3255 adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3256 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3257 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3258 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3259 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3260 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3261 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3262 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3263 VSS col_n[2] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3264 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3265 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3266 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3267 VSS col_n[6] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3268 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3269 adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3270 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3271 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3272 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3273 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3274 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3275 vcom VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3276 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3277 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3278 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vint2 en_n_bit[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3279 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3280 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3281 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3282 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3283 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3284 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3285 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3286 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3287 VDD sample adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3288 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3289 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3290 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3291 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vint2 en_n_bit[1] adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3292 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3293 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3294 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3295 VSS col_n[10] adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3296 VDD sample_n adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3297 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3298 VSS col_n[0] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3299 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3300 VSS col_n[11] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3301 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3302 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3303 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3304 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3305 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3306 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3307 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3308 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3309 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3310 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3311 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3312 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3313 VSS VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3314 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3315 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3316 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3317 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3318 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3319 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3320 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3321 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3322 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3323 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3324 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3325 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3326 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3327 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3328 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3329 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3330 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3331 VSS col_n[7] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3332 adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3333 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3334 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3335 VSS col_n[1] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3336 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3337 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3338 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3339 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3340 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3341 vcom VSS adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3342 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3343 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3344 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3345 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3346 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3347 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3348 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3349 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3350 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3351 adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3352 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3353 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3354 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3355 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3356 VSS col_n[5] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3357 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3358 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3359 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3360 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3361 VSS col_n[8] adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3362 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3363 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3364 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3365 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3366 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3367 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3368 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3369 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3370 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3371 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3372 VSS col_n[12] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3373 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3374 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3375 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X3376 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3377 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3378 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3379 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3380 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3381 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3382 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3383 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3384 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3385 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3386 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3387 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3388 VSS col_n[9] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3389 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3390 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3391 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3392 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3393 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3394 VSS col_n[3] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3395 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3396 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3397 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3398 VSS VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3399 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3400 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3401 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3402 VSS VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3403 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3404 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3405 VSS col_n[15] adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3406 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3407 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3408 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3409 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3410 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3411 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3412 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3413 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3414 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3415 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3416 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3417 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3418 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3419 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3420 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3421 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3422 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3423 VSS sample adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3424 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3425 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3426 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3427 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3428 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3429 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3430 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3431 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3432 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3433 VSS VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3434 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3435 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3436 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3437 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3438 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3439 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3440 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3441 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3442 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3443 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3444 VSS col_n[13] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3445 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3446 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3447 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3448 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3449 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3450 adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3451 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3452 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3453 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3454 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3455 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3456 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3457 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3458 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3459 ctop sw analog_in VSS sky130_fd_pr__nfet_01v8 ad=1.45e+11p pd=1.58e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=500000u
X3460 VDD VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3461 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3462 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3463 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3464 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3465 VSS col_n[11] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3466 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3467 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3468 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3469 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3470 VSS col_n[11] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3471 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3472 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3473 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3474 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3475 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3476 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3477 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3478 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3479 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3480 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3481 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3482 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3483 VSS col_n[3] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3484 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3485 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3486 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3487 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3488 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3489 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3490 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3491 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3492 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3493 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3494 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3495 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3496 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3497 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3498 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3499 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3500 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3501 VSS col_n[14] adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3502 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3503 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3504 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3505 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X3506 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3507 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3508 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3509 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3510 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3511 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3512 VDD VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3513 VSS col_n[7] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3514 VSS col_n[3] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3515 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3516 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3517 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3518 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3519 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3520 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3521 VSS VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3522 VDD colon_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3523 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3524 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3525 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3526 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3527 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3528 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3529 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3530 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3531 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3532 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3533 VDD colon_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3534 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3535 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3536 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3537 VSS col_n[12] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3538 VSS col_n[5] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3539 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3540 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3541 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3542 VSS col_n[8] adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3543 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3544 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3545 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3546 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3547 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3548 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3549 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3550 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3551 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3552 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3553 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3554 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3555 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3556 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3557 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X3558 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3559 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3560 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3561 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3562 VSS col_n[3] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3563 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3564 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3565 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3566 VDD sample_n adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3567 VSS col_n[14] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3568 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3569 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3570 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3571 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3572 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3573 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3574 adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3575 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3576 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3577 vcom VSS adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3578 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3579 adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3580 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3581 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3582 vcom VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3583 VDD VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3584 vcom VSS adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3585 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3586 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3587 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3588 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3589 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3590 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3591 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3592 VSS col_n[10] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3593 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3594 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3595 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3596 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3597 VSS col_n[0] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3598 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3599 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3600 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3601 VSS col_n[4] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3602 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3603 adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3604 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3605 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3606 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3607 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3608 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3609 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3610 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3611 VSS VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3612 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3613 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3614 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3615 adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3616 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3617 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3618 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3619 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3620 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3621 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3622 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3623 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3624 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3625 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3626 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3627 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3628 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3629 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3630 vcom VSS adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3631 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3632 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3633 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3634 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3635 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3636 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3637 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3638 VSS col_n[15] adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3639 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3640 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3641 vcom VSS adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3642 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3643 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3644 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3645 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3646 VSS col_n[1] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3647 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3648 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3649 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3650 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3651 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3652 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3653 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3654 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3655 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3656 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3657 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3658 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3659 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3660 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3661 adc_array_wafflecap_8_Dummy_0[8]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3662 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3663 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3664 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3665 VSS col_n[5] adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3666 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3667 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3668 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3669 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3670 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3671 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3672 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3673 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3674 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3675 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3676 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3677 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3678 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3679 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3680 adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3681 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3682 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3683 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3684 VSS col_n[9] adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3685 VDD en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3686 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3687 VSS col_n[3] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3688 VSS col_n[7] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3689 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3690 VSS sample_n adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3691 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3692 VSS VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3693 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3694 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3695 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3696 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3697 VSS col_n[11] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3698 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3699 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3700 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3701 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3702 VSS col_n[6] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3703 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3704 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3705 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3706 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3707 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3708 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3709 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3710 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3711 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3712 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3713 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3714 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3715 VSS col_n[8] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3716 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3717 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3718 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3719 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3720 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3721 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3722 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3723 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3724 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3725 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3726 VSS col_n[14] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3727 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3728 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3729 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3730 VSS col_n[14] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3731 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3732 VSS col_n[13] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3733 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3734 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3735 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3736 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3737 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3738 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3739 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3740 VDD VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3741 VDD VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3742 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3743 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3744 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3745 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3746 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3747 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3748 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3749 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3750 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3751 VSS sample adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3752 VSS col_n[9] adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3753 adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3754 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3755 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3756 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3757 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3758 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3759 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3760 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3761 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3762 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3763 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3764 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3765 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3766 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3767 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3768 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3769 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3770 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3771 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3772 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3773 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3774 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3775 adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3776 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3777 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3778 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3779 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3780 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3781 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3782 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3783 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3784 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3785 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3786 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3787 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3788 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3789 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3790 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3791 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3792 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3793 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3794 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3795 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3796 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3797 VDD VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3798 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3799 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3800 VSS col_n[15] adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3801 VSS col_n[15] adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3802 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3803 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3804 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3805 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3806 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3807 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3808 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3809 VSS col_n[7] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3810 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3811 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3812 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3813 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3814 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3815 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3816 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3817 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3818 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3819 VSS col_n[1] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3820 VSS col_n[10] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3821 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3822 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3823 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3824 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3825 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3826 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3827 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3828 VSS col_n[12] adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3829 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3830 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3831 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3832 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3833 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3834 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3835 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3836 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3837 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3838 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3839 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3840 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3841 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3842 VSS col_n[5] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3843 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3844 VDD sample adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3845 VSS col_n[8] adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3846 adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_Dummy_5[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3847 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint1 en_n_bit[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3848 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3849 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3850 analog_in sw ctop VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=500000u l=500000u
X3851 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3852 vcom VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3853 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3854 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3855 VSS col_n[14] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3856 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3857 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3858 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3859 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3860 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3861 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3862 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3863 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3864 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3865 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3866 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3867 VSS col_n[7] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3868 VSS col_n[3] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3869 VDD VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3870 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3871 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3872 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3873 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3874 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3875 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3876 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3877 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3878 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3879 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3880 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3881 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3882 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3883 VSS col_n[6] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3884 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3885 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3886 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3887 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3888 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3889 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3890 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3891 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3892 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3893 VSS sample_n adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3894 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3895 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3896 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3897 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3898 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X3899 VSS col_n[1] adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3900 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3901 VSS col_n[12] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3902 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3903 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3904 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3905 adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3906 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X3907 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3908 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3909 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3910 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3911 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3912 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3913 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3914 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3915 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3916 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3917 VSS col_n[9] adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3918 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3919 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3920 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3921 VSS col_n[9] adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3922 adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3923 adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3924 VSS col_n[15] adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3925 adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3926 vcom VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3927 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3928 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3929 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3930 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3931 VSS VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3932 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3933 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3934 VSS col_n[2] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3935 VSS VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3936 VSS col_n[8] adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3937 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3938 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3939 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3940 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3941 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3942 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3943 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3944 vcom VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3945 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3946 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3947 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3948 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3949 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3950 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3951 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3952 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3953 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3954 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X3955 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3956 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3957 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3958 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3959 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3960 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3961 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3962 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3963 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3964 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3965 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3966 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3967 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3968 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3969 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3970 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3971 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X3972 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3973 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3974 VSS col_n[13] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3975 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3976 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3977 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3978 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3979 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X3980 adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3981 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3982 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3983 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3984 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3985 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X3986 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3987 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3988 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X3989 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3990 VSS col_n[10] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3991 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3992 VSS col_n[10] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3993 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3994 VSS col_n[11] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3995 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X3996 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X3997 VSS col_n[11] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3998 adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3999 VSS col_n[3] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4000 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4001 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4002 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4003 VSS col_n[7] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4004 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4005 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4006 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint2 en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4007 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4008 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4009 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4010 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4011 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4012 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4013 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4014 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4015 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4016 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4017 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4018 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4019 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4020 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4021 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4022 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4023 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4024 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4025 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4026 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4027 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4028 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4029 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4030 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4031 VSS col_n[5] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4032 VSS col_n[8] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4033 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4034 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4035 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4036 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4037 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4038 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4039 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4040 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4041 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4042 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4043 VSS col_n[4] adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4044 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4045 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4046 VDD VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4047 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4048 VSS col_n[9] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4049 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4050 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4051 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4052 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4053 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4054 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4055 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4056 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4057 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4058 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4059 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4060 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4061 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4062 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4063 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4064 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4065 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4066 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4067 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4068 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4069 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4070 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4071 VSS col_n[12] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4072 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4073 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4074 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4075 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4076 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4077 VSS col_n[12] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4078 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4079 adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4080 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4081 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4082 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4083 adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4084 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4085 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4086 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4087 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4088 VSS sample adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4089 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4090 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4091 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X4092 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4093 VSS sample_n adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4094 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4095 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4096 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4097 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4098 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint2 en_n_bit[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4099 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4100 VSS sample adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4101 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4102 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4103 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4104 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4105 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4106 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4107 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X4108 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4109 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4110 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4111 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4112 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4113 VSS col_n[15] adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4114 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4115 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4116 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4117 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4118 vcom VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4119 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4120 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4121 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4122 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4123 VSS col_n[10] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4124 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4125 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4126 adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4127 VSS col_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4128 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4129 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4130 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4131 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4132 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4133 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4134 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4135 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4136 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4137 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4138 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4139 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4140 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4141 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4142 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4143 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4144 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4145 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4146 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4147 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4148 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4149 VSS col_n[13] adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4150 VSS col_n[13] adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4151 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4152 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4153 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4154 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4155 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4156 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4157 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4158 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4159 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4160 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4161 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4162 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4163 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4164 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4165 adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4166 VSS col_n[5] adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4167 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4168 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4169 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4170 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4171 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4172 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4173 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4174 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4175 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4176 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4177 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4178 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4179 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4180 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4181 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4182 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4183 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4184 VSS en_n_bit[2] adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4185 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4186 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4187 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4188 vcom VSS adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4189 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4190 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4191 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4192 VSS col_n[15] adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4193 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4194 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4195 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4196 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4197 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4198 VSS col_n[7] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4199 VSS col_n[3] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4200 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4201 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4202 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4203 VDD sample adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4204 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4205 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4206 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4207 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4208 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4209 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4210 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4211 VSS col_n[12] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4212 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4213 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4214 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4215 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4216 VSS col_n[6] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4217 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint1 row_n[21] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4218 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4219 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4220 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4221 adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4222 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4223 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4224 VSS col_n[5] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4225 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4226 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4227 VSS col_n[8] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4228 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4229 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4230 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4231 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4232 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4233 adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4234 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4235 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4236 VSS col_n[1] adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4237 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4238 VSS col_n[4] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4239 vcom VSS adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4240 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4241 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4242 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4243 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4244 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4245 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4246 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4247 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4248 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4249 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4250 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4251 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4252 VSS sample_n adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4253 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4254 adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4255 adc_array_wafflecap_8_Dummy_0[6]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4256 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4257 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4258 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4259 VSS col_n[11] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4260 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4261 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4262 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4263 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4264 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4265 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4266 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4267 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4268 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4269 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4270 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4271 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4272 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4273 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4274 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4275 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4276 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4277 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4278 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4279 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4280 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4281 VSS col_n[13] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4282 adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4283 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4284 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4285 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4286 VDD VSS adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4287 VSS col_n[0] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4288 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4289 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4290 VSS col_n[14] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4291 VSS sample adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4292 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4293 VSS col_n[14] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4294 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4295 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4296 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4297 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4298 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4299 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4300 adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4301 VSS VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4302 VDD VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4303 adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4304 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4305 VDD VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4306 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4307 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4308 adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4309 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4310 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4311 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4312 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4313 adc_array_wafflecap_8_8_0[8|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4314 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4315 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4316 VSS col_n[10] adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4317 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4318 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4319 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4320 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4321 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4322 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4323 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4324 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4325 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4326 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4327 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4328 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4329 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4330 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4331 adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4332 adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4333 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4334 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4335 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4336 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4337 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4338 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4339 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4340 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4341 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4342 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4343 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4344 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4345 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4346 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4347 adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4348 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4349 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4350 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4351 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4352 vcom VSS adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4353 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4354 vcom VSS adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4355 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4356 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=7.44e+11p pd=6.66e+06u as=0p ps=0u w=800000u l=150000u
X4357 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4358 adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4359 VSS col_n[5] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4360 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4361 VSS col_n[15] adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4362 VSS col_n[15] adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4363 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4364 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4365 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4366 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4367 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4368 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4369 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4370 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4371 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4372 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4373 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4374 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4375 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4376 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4377 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4378 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4379 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4380 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4381 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4382 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4383 VSS col_n[3] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4384 VSS col_n[10] adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4385 adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4386 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4387 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4388 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4389 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4390 adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4391 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4392 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4393 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4394 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4395 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4396 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4397 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4398 VSS col_n[6] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4399 VSS col_n[2] adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4400 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4401 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4402 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4403 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4404 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4405 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4406 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4407 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4408 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4409 VSS col_n[8] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4410 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4411 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4412 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4413 VSS col_n[15] adc_array_wafflecap_8_8_0[15|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4414 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4415 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4416 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4417 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4418 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4419 VSS col_n[1] adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4420 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4421 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4422 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4423 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4424 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4425 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4426 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4427 adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4428 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4429 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4430 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4431 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4432 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4433 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4434 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4435 adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4436 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4437 VSS sample adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4438 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4439 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4440 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4441 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4442 VSS col_n[8] adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4443 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4444 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4445 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4446 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4447 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4448 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4449 adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4450 vcom VSS adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4451 adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4452 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4453 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4454 VSS col_n[13] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4455 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4456 adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4457 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4458 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4459 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4460 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4461 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4462 adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4463 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4464 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4465 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4466 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4467 adc_array_wafflecap_8_Dummy_3[3]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4468 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4469 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4470 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4471 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4472 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4473 VSS col_n[9] adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4474 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4475 VSS col_n[9] adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4476 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4477 VSS col_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4478 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4479 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4480 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4481 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4482 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4483 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4484 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4485 adc_array_wafflecap_8_8_0[8|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4486 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4487 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4488 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4489 VSS VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4490 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4491 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4492 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4493 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4494 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4495 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4496 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4497 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4498 adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4499 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4500 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4501 VSS col_n[7] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4502 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4503 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4504 VSS col_n[3] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4505 adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4506 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4507 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4508 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X4509 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4510 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4511 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4512 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4513 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4514 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4515 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4516 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4517 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4518 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4519 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4520 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4521 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4522 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4523 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4524 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4525 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4526 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4527 adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4528 vcom VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4529 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4530 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4531 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4532 VSS VSS adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X4533 VSS col_n[13] adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4534 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4535 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4536 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4537 VSS col_n[5] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4538 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4539 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4540 VDD sample adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4541 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4542 VSS VDD adc_array_wafflecap_8_Dummy_4[27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4543 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4544 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4545 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4546 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4547 adc_array_wafflecap_8_8_0[12|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4548 VSS col_n[10] adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4549 VSS col_n[10] adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4550 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4551 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4552 VSS col_n[4] adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4553 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4554 VSS col_n[11] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4555 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4556 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4557 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4558 adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4559 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4560 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4561 VSS col_n[3] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4562 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4563 adc_array_wafflecap_8_8_0[9|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4564 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4565 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4566 adc_array_wafflecap_8_8_0[9|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4567 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4568 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4569 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4570 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4571 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4572 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4573 adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4574 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4575 adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4576 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4577 VSS sample_n adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4578 adc_array_wafflecap_8_Dummy_4[16]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4579 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4580 VSS col_n[6] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4581 VSS col_n[2] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4582 adc_array_wafflecap_8_Dummy_4[6]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4583 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4584 adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4585 adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4586 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4587 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4588 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4589 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4590 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4591 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4592 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4593 vcom VSS adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4594 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4595 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4596 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4597 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4598 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4599 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4600 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4601 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4602 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4603 VSS col_n[1] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4604 VSS col_n[10] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4605 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4606 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4607 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4608 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4609 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4610 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4611 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.44e+11p ps=6.66e+06u w=800000u l=150000u
X4612 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4613 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4614 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.604e+11p ps=2.92e+06u w=420000u l=150000u
X4615 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4616 adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4617 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4618 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4619 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4620 adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4621 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4622 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4623 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4624 adc_array_wafflecap_8_8_0[5|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4625 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4626 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4627 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4628 adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4629 VSS col_n[12] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4630 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4631 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4632 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4633 VSS col_n[12] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4634 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4635 VSS col_n[8] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4636 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4637 adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4638 adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4639 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4640 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4641 adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4642 adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4643 adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4644 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4645 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4646 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4647 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4648 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4649 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4650 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4651 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4652 adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4653 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4654 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4655 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4656 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4657 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4658 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4659 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4660 vcom VSS adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4661 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4662 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4663 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4664 adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4665 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4666 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4667 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4668 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4669 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4670 adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4671 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4672 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4673 adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4674 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4675 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4676 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4677 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4678 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4679 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4680 VSS col_n[10] adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4681 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4682 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4683 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4684 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4685 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint1 VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4686 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4687 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4688 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4689 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4690 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4691 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4692 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4693 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4694 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4695 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4696 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4697 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4698 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4699 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4700 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4701 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4702 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4703 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4704 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4705 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4706 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4707 VSS col_n[3] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4708 VSS col_n[13] adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4709 VSS col_n[13] adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4710 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4711 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4712 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4713 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4714 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4715 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4716 adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4717 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4718 VSS VDD adc_array_wafflecap_8_Dummy_4[12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4719 adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4720 VSS VDD adc_array_wafflecap_8_Dummy_4[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4721 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4722 adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4723 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4724 vcom VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4725 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4726 adc_array_wafflecap_8_8_0[12|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4727 adc_array_wafflecap_8_8_0[12|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4728 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4729 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4730 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4731 VSS col_n[8] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4732 adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4733 adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4734 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4735 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4736 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4737 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4738 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4739 vcom VSS adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4740 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4741 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4742 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4743 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4744 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4745 VSS col_n[1] adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4746 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4747 VSS col_n[4] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4748 VSS col_n[0] adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4749 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4750 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4751 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4752 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4753 adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4754 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4755 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4756 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4757 adc_array_wafflecap_8_8_0[15|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4758 VSS col_n[13] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4759 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4760 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4761 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4762 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4763 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4764 adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4765 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4766 VSS col_n[8] adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4767 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4768 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4769 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4770 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4771 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4772 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4773 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4774 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4775 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4776 adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4777 adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4778 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4779 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4780 adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4781 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4782 adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4783 adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4784 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4785 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4786 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4787 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4788 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4789 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4790 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4791 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4792 adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4793 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4794 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4795 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4796 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4797 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4798 adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4799 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4800 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4801 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4802 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4803 adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4804 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X4805 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4806 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4807 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4808 adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4809 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4810 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4811 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4812 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4813 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4814 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4815 vcom VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X4816 adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4817 adc_array_wafflecap_8_8_0[8|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4818 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4819 VSS col_n[8] adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4820 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4821 adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4822 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4823 VDD sample_n adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4824 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4825 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4826 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4827 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4828 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4829 VSS col_n[1] adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4830 adc_array_wafflecap_8_8_0[15|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4831 VSS col_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4832 adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4833 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4834 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4835 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4836 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4837 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4838 adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4839 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4840 VSS col_n[14] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4841 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4842 adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4843 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4844 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4845 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4846 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4847 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4848 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4849 adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4850 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4851 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4852 adc_array_wafflecap_8_8_0[3|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4853 adc_array_wafflecap_8_Dummy_0[4]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4854 adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4855 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4856 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4857 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4858 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4859 VDD VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4860 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4861 VSS col_n[5] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4862 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4863 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4864 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4865 adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4866 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4867 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4868 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4869 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4870 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4871 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4872 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4873 adc_array_wafflecap_8_8_0[1|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4874 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4875 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4876 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4877 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4878 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4879 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4880 VDD VSS adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4881 adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4882 adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4883 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4884 VDD sample_n adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4885 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4886 VSS col_n[3] adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4887 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4888 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4889 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4890 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4891 VDD sample adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4892 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4893 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4894 VSS col_n[14] adc_array_wafflecap_8_8_0[14|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4895 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4896 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4897 adc_array_wafflecap_8_8_0[11|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4898 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4899 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4900 vcom VSS adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4901 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4902 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4903 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4904 VSS col_n[6] adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4905 VSS col_n[2] adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4906 VDD VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4907 vcom VSS adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4908 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4909 adc_array_wafflecap_8_8_0[8|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4910 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4911 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4912 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4913 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4914 adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4915 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4916 adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4917 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4918 adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4919 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4920 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4921 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4922 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4923 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4924 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4925 adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4926 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4927 adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4928 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4929 VSS col_n[1] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4930 adc_array_wafflecap_8_8_0[14|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4931 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4932 VSS col_n[4] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4933 VSS col_n[0] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4934 adc_array_wafflecap_8_8_0[14|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4935 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4936 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4937 adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4938 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4939 adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4940 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4941 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4942 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4943 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4944 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4945 adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4946 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4947 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4948 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4949 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4950 adc_array_wafflecap_8_8_0[3|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4951 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4952 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4953 adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4954 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X4955 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4956 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4957 VSS col_n[8] adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4958 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4959 adc_array_wafflecap_8_8_0[10|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4960 adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4961 adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4962 adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4963 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4964 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4965 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4966 VSS VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4967 adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4968 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4969 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4970 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4971 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4972 VSS col_n[15] adc_array_wafflecap_8_8_0[15|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4973 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4974 adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4975 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4976 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4977 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4978 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4979 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4980 adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4981 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4982 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4983 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4984 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4985 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4986 adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4987 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4988 adc_array_wafflecap_8_8_0[3|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4989 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X4990 adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4991 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4992 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4993 adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4994 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4995 adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4996 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4997 adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X4998 adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X4999 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5000 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5001 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5002 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5003 adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5004 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5005 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5006 adc_array_wafflecap_8_8_0[15|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5007 adc_array_wafflecap_8_8_0[15|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5008 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5009 adc_array_wafflecap_8_8_0[6|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5010 adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5011 adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5012 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5013 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5014 adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5015 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5016 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5017 adc_array_wafflecap_8_8_0[4|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5018 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint2 row_n[22] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5019 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5020 VSS sample adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5021 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5022 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5023 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5024 VSS col_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5025 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5026 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5027 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5028 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5029 adc_array_wafflecap_8_8_0[10|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5030 adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5031 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5032 VSS col_n[11] adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5033 adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5034 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5035 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5036 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5037 vcom VSS adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5038 VSS col_n[9] adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5039 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5040 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5041 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5042 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5043 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5044 adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5045 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5046 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5047 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5048 VDD sample_n adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5049 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5050 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5051 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5052 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5053 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5054 adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5055 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5056 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5057 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5058 adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5059 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5060 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5061 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5062 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5063 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5064 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5065 VSS col_n[14] adc_array_wafflecap_8_8_0[14|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5066 adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5067 VSS col_n[14] adc_array_wafflecap_8_8_0[14|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5068 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5069 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5070 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5071 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5072 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5073 VDD VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5074 VDD sample adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5075 adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5076 VSS VSS adc_array_wafflecap_8_Dummy_1[6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5077 VDD VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5078 adc_array_wafflecap_8_8_0[7|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5079 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5080 adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5081 adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5082 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5083 adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5084 adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5085 adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5086 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5087 adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5088 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5089 VSS col_n[9] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5090 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5091 VSS col_n[2] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5092 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5093 VSS col_n[6] adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5094 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5095 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5096 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5097 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5098 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5099 adc_array_wafflecap_8_8_0[6|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5100 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5101 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5102 adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5103 VSS col_n[11] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5104 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5105 VDD VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5106 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5107 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5108 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5109 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5110 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5111 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5112 adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5113 adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5114 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5115 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5116 VSS col_n[1] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5117 adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5118 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5119 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5120 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5121 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5122 adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_Dummy_5[7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5123 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5124 adc_array_wafflecap_8_8_0[9|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5125 adc_array_wafflecap_8_8_0[9|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5126 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5127 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5128 adc_array_wafflecap_8_8_0[5|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5129 adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5130 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5131 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5132 adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5133 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5134 adc_array_wafflecap_8_Dummy_5[15]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5135 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5136 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5137 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5138 VSS VSS adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.688e+11p ps=2.96e+06u w=420000u l=150000u
X5139 VSS col_n[15] adc_array_wafflecap_8_8_0[15|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5140 VSS col_n[8] adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5141 adc_array_wafflecap_8_Dummy_4[9]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5142 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5143 adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5144 adc_array_wafflecap_8_Dummy_1[3]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5145 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5146 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5147 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5148 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5149 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5150 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5151 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5152 adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5153 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5154 VSS col_n[10] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5155 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5156 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5157 adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5158 adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5159 adc_array_wafflecap_8_8_0[3|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5160 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5161 adc_array_wafflecap_8_Dummy_2[1]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5162 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5163 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5164 adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5165 VSS col_n[6] adc_array_wafflecap_8_8_0[6|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5166 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5167 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5168 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5169 adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5170 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5171 VDD VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5172 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5173 adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5174 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5175 adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5176 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5177 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5178 adc_array_wafflecap_8_8_0[5|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5179 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5180 adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5181 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5182 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5183 VSS col_n[12] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5184 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5185 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5186 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5187 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5188 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5189 adc_array_wafflecap_8_8_0[10|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5190 adc_array_wafflecap_8_8_0[10|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5191 adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5192 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5193 adc_array_wafflecap_8_8_0[1|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5194 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5195 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5196 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5197 VSS col_n[7] adc_array_wafflecap_8_8_0[7|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5198 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5199 adc_array_wafflecap_8_8_0[0|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5200 VSS col_n[3] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5201 adc_array_wafflecap_8_8_0[11|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5202 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5203 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5204 adc_array_wafflecap_8_8_0[4|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5205 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5206 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5207 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5208 adc_array_wafflecap_8_8_0[3|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5209 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5210 adc_array_wafflecap_8_8_0[6|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5211 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5212 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5213 adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5214 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5215 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint1 row_n[16] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5216 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5217 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5218 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5219 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5220 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5221 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5222 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5223 VDD sample adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5224 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5225 adc_array_wafflecap_8_8_0[2|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5226 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5227 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5228 VDD sample_n adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5229 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5230 adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5231 adc_array_wafflecap_8_8_0[4|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5232 VDD sample adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5233 adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5234 adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5235 VSS col_n[12] adc_array_wafflecap_8_8_0[12|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5236 adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5237 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5238 adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5239 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5240 adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5241 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5242 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5243 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5244 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5245 adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5246 VSS col_n[4] adc_array_wafflecap_8_8_0[4|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5247 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5248 VSS col_n[0] adc_array_wafflecap_8_8_0[0|10]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5249 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5250 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5251 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5252 VSS col_n[9] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5253 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5254 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5255 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5256 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5257 adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5258 VSS col_n[9] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5259 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5260 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5261 adc_array_wafflecap_8_8_0[7|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5262 adc_array_wafflecap_8_8_0[6|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5263 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5264 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5265 adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5266 adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5267 VSS VDD adc_array_wafflecap_8_Dummy_4[15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5268 adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5269 adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5270 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5271 VSS VDD adc_array_wafflecap_8_Dummy_4[5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5272 VSS col_n[8] adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5273 adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5274 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5275 adc_array_wafflecap_8_8_0[12|15]/adc_array_circuit_150n_0/vint2 row_n[15] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5276 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5277 VSS col_n[2] adc_array_wafflecap_8_8_0[2|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5278 adc_array_wafflecap_8_8_0[12|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5279 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5280 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5281 adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5282 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5283 VSS col_n[11] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5284 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5285 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5286 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5287 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5288 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5289 adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5290 adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5291 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5292 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5293 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5294 adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5295 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5296 adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|5]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5297 adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|15]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5298 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5299 adc_array_wafflecap_8_8_0[8|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5300 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5301 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5302 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5303 adc_array_wafflecap_8_Dummy_5[4]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5304 vcom VSS adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5305 VSS col_n[1] adc_array_wafflecap_8_8_0[1|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5306 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5307 adc_array_wafflecap_8_Dummy_0[5]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5308 adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5309 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5310 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5311 VSS col_n[14] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5312 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5313 VSS col_n[13] adc_array_wafflecap_8_8_0[13|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5314 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5315 adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5316 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5317 VDD VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5318 adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5319 adc_array_wafflecap_8_8_0[14|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5320 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5321 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5322 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5323 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5324 adc_array_wafflecap_8_Dummy_5[10]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5325 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5326 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5327 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5328 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5329 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5330 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5331 adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5332 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5333 VSS col_n[10] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5334 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5335 adc_array_wafflecap_8_8_0[1|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5336 adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5337 adc_array_wafflecap_8_Dummy_6/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5338 VSS col_n[1] adc_array_wafflecap_8_8_0[1|28]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5339 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5340 adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5341 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5342 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5343 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5344 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5345 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5346 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5347 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5348 adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5349 adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5350 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5351 adc_array_wafflecap_8_8_0[13|3]/adc_array_circuit_150n_0/vint2 row_n[3] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5352 adc_array_wafflecap_8_8_0[13|13]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5353 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5354 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5355 adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5356 adc_array_wafflecap_8_8_0[3|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5357 adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5358 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5359 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5360 VSS VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5361 adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5362 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5363 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5364 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5365 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vint1 row_n[12] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5366 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5367 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5368 adc_array_wafflecap_8_8_0[2|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5369 VSS sample adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5370 adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5371 adc_array_wafflecap_8_8_0[2|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5372 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5373 adc_array_wafflecap_8_8_0[5|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5374 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5375 adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5376 adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5377 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5378 adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_4_0/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5379 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.64e+07u l=1.6e+07u
X5380 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5381 adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5382 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5383 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5384 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5385 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5386 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5387 adc_array_wafflecap_8_8_0[1|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5388 adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5389 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5390 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5391 adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5392 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5393 adc_array_wafflecap_8_8_0[0|5]/adc_array_circuit_150n_0/vint2 row_n[5] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5394 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5395 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5396 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5397 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5398 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5399 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5400 adc_array_wafflecap_8_8_0[6|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5401 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5402 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vint1 row_n[2] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5403 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5404 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5405 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5406 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5407 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5408 adc_array_wafflecap_8_8_0[8|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5409 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5410 VSS col_n[12] adc_array_wafflecap_8_8_0[12|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5411 adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5412 adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5413 VSS col_n[12] adc_array_wafflecap_8_8_0[12|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5414 adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5415 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5416 vcom VSS adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.386e+11p ps=1.5e+06u w=420000u l=150000u
X5417 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5418 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5419 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5420 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5421 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5422 VDD sample adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5423 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5424 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5425 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5426 adc_array_wafflecap_8_8_0[4|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5427 adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5428 adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/vint1 row_n[1] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5429 adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5430 adc_array_wafflecap_8_8_0[7|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5431 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5432 adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5433 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5434 adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5435 adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5436 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5437 VSS col_n[0] adc_array_wafflecap_8_8_0[0|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5438 adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5439 VSS col_n[4] adc_array_wafflecap_8_8_0[4|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5440 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5441 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5442 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5443 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5444 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5445 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5446 VSS col_n[15] adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5447 adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5448 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5449 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5450 adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5451 adc_array_wafflecap_8_Dummy_4[22]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5452 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5453 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5454 adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5455 adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5456 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5457 adc_array_wafflecap_8_8_0[2|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5458 adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5459 vcom VSS adc_array_wafflecap_8_Dummy_4[17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5460 VSS col_n[8] adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5461 VDD VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5462 VDD VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5463 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5464 vcom VSS adc_array_wafflecap_8_Dummy_4[7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5465 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5466 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5467 adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5468 adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5469 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5470 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5471 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5472 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5473 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5474 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5475 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5476 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5477 adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5478 adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5479 adc_array_wafflecap_8_8_0[8|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5480 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5481 VDD colon_n[8] adc_array_wafflecap_8_Dummy_5[8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5482 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5483 VDD VSS adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5484 VSS col_n[13] adc_array_wafflecap_8_8_0[13|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5485 adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5486 adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5487 adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5488 adc_array_wafflecap_8_8_0[14|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5489 adc_array_wafflecap_8_8_0[3|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5490 adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5491 adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vint1 row_n[31] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5492 adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5493 adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_2[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5494 adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5495 adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5496 adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5497 VSS col_n[6] adc_array_wafflecap_8_8_0[6|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5498 adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5499 adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5500 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5501 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5502 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5503 adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5504 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5505 adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5506 adc_array_wafflecap_8_8_0[14|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5507 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5508 VSS col_n[9] adc_array_wafflecap_8_8_0[9|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5509 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5510 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5511 adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5512 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5513 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5514 adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5515 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5516 VSS VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5517 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5518 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5519 VSS col_n[4] adc_array_wafflecap_8_8_0[4|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5520 VSS col_n[15] adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5521 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5522 adc_array_wafflecap_8_2_0/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5523 adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5524 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|15]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5525 adc_array_wafflecap_8_8_0[4|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5526 VSS col_n[1] adc_array_wafflecap_8_8_0[1|29]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5527 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5528 adc_array_wafflecap_8_Dummy_4[33]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5529 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|5]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5530 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5531 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5532 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5533 adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5534 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5535 adc_array_wafflecap_8_8_0[3|10]/adc_array_circuit_150n_0/vint2 row_n[10] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5536 adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5537 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5538 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5539 adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5540 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5541 adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5542 adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5543 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5544 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5545 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5546 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5547 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5548 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5549 VSS col_n[5] adc_array_wafflecap_8_8_0[5|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5550 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5551 adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5552 adc_array_wafflecap_8_8_0[2|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5553 adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5554 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5555 adc_array_wafflecap_8_8_0[15|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5556 adc_array_wafflecap_8_8_0[4|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5557 adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5558 adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5559 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5560 adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5561 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5562 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5563 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5564 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5565 adc_array_wafflecap_8_8_0[0|7]/adc_array_circuit_150n_0/vint2 row_n[7] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5566 adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5567 adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5568 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5569 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5570 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5571 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5572 VSS col_n[11] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5573 adc_array_wafflecap_8_8_0[6|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5574 adc_array_wafflecap_8_8_0[2|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5575 adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5576 adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_1_0/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5577 adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5578 adc_array_wafflecap_8_8_0[11|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5579 adc_array_wafflecap_8_8_0[11|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5580 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint2 row_n[14] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5581 adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5582 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5583 adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint2 row_n[13] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5584 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5585 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5586 adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5587 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5588 VSS col_n[2] adc_array_wafflecap_8_8_0[2|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5589 adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5590 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5591 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5592 adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n sample VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5593 adc_array_wafflecap_8_8_0[9|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5594 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5595 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5596 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5597 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5598 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5599 adc_array_wafflecap_8_Dummy_4[21]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5600 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5601 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5602 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5603 adc_array_wafflecap_8_8_0[4|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5604 adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5605 adc_array_wafflecap_8_8_0[7|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5606 adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5607 VSS col_n[14] adc_array_wafflecap_8_8_0[14|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5608 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5609 adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|9]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5610 adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5611 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint1 row_n[9] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5612 VSS col_n[14] adc_array_wafflecap_8_8_0[14|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5613 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5614 adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5615 VSS col_n[1] adc_array_wafflecap_8_8_0[1|1]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5616 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5617 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5618 VSS col_n[0] adc_array_wafflecap_8_8_0[0|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5619 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5620 VDD VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5621 adc_array_wafflecap_8_8_0[13|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5622 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5623 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5624 VDD VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5625 adc_array_wafflecap_8_8_0[13|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5626 adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5627 adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5628 adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|11]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5629 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5630 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5631 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5632 adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|22]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5633 adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5634 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5635 adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5636 VSS col_n[10] adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5637 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5638 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5639 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5640 VSS col_n[8] adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5641 adc_array_wafflecap_8_Dummy_5[2]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5642 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5643 adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5644 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5645 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5646 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vint2 colon_n[15] adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5647 VSS col_n[12] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5648 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5649 VSS col_n[1] adc_array_wafflecap_8_8_0[1|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5650 adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|21]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5651 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5652 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5653 adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5654 adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5655 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5656 VSS col_n[7] adc_array_wafflecap_8_8_0[7|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5657 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5658 adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5659 adc_array_wafflecap_8_8_0[8|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5660 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5661 adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5662 adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5663 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5664 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5665 VDD colon_n[13] adc_array_wafflecap_8_Dummy_5[13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5666 adc_array_wafflecap_8_8_0[3|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5667 adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5668 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5669 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5670 adc_array_wafflecap_8_8_0[10|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5671 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5672 adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5673 VSS VSS adc_array_wafflecap_8_Dummy_1[4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5674 VDD colon_n[3] adc_array_wafflecap_8_Dummy_5[3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5675 adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5676 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5677 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5678 adc_array_wafflecap_8_8_0[9|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5679 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint1 row_n[13] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5680 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5681 VSS col_n[6] adc_array_wafflecap_8_8_0[6|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5682 adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5683 VSS col_n[15] adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5684 VSS col_n[15] adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5685 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5686 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint1 row_n[27] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5687 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vdrv col_n[1] adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5688 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv col_n[14] adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5689 adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5690 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5691 adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5692 adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5693 adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5694 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5695 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=2.64e+11p pd=2.26e+06u as=0p ps=0u w=800000u l=150000u
X5696 adc_array_wafflecap_8_8_0[1|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5697 adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5698 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5699 adc_array_wafflecap_8_8_0[0|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5700 adc_array_wafflecap_8_8_0[0|0]/adc_array_circuit_150n_0/vint2 row_n[0] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5701 VSS col_n[1] adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5702 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5703 VSS col_n[10] adc_array_wafflecap_8_8_0[10|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5704 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5705 VDD sample_n adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5706 adc_array_wafflecap_8_8_0[3|12]/adc_array_circuit_150n_0/vint2 row_n[12] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5707 adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5708 adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5709 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5710 adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_4[32]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5711 adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5712 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5713 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5714 vcom adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[12]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5715 adc_array_wafflecap_8_8_0[8|23]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5716 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5717 adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5718 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5719 adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/cbot VDD adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5720 adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5721 adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5722 VSS VSS adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5723 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5724 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5725 adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5726 adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5727 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5728 adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5729 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5730 adc_array_wafflecap_8_Dummy_1[1]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5731 adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5732 adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5733 adc_array_wafflecap_8_8_0[11|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5734 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5735 adc_array_wafflecap_8_8_0[4|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5736 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5737 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5738 adc_array_wafflecap_8_8_0[10|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5739 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5740 adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5741 adc_array_wafflecap_8_8_0[13|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5742 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5743 adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|30]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5744 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5745 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5746 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5747 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5748 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5749 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5750 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5751 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5752 adc_array_wafflecap_8_8_0[9|28]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5753 adc_array_wafflecap_8_8_0[6|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5754 adc_array_wafflecap_8_8_0[2|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5755 adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5756 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|24]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5757 VSS col_n[8] adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5758 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample sample_n VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5759 adc_array_wafflecap_8_8_0[5|4]/adc_array_circuit_150n_0/vint2 row_n[4] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5760 adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5761 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5762 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5763 VDD VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5764 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5765 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5766 VSS col_n[2] adc_array_wafflecap_8_8_0[2|11]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5767 adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5768 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5769 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5770 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=2.688e+11p pd=2.96e+06u as=0p ps=0u w=420000u l=150000u
X5771 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5772 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5773 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5774 adc_array_wafflecap_8_8_0[8|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5775 VSS col_n[13] adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5776 adc_array_wafflecap_8_8_0[12|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5777 adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5778 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5779 adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5780 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5781 adc_array_wafflecap_8_8_0[7|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5782 VDD VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5783 adc_array_wafflecap_8_8_0[1|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5784 adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[18]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5785 adc_array_wafflecap_8_8_0[14|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5786 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5787 adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|11]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5788 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vint1 row_n[11] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5789 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5790 adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5791 adc_array_wafflecap_8_8_0[0|30]/adc_array_circuit_150n_0/vint2 row_n[30] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5792 adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vint2 colon_n[0] adc_array_wafflecap_8_8_0[0|18]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5793 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5794 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5795 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|28]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5796 vcom adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5797 adc_array_wafflecap_8_8_0[11|25]/adc_array_circuit_150n_0/vint1 row_n[25] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5798 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5799 VSS col_n[9] adc_array_wafflecap_8_8_0[9|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5800 adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_0[3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5801 VSS col_n[9] adc_array_wafflecap_8_8_0[9|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5802 adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5803 VSS col_n[15] adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5804 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5805 adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5806 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5807 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5808 adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5809 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5810 VSS VDD adc_array_wafflecap_8_Dummy_4[8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5811 VDD colon_n[6] adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5812 adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vdrv VDD adc_array_wafflecap_8_Dummy_4[24]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5813 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5814 VSS col_n[8] adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5815 VDD VSS sky130_fd_pr__cap_mim_m3_1 l=1.72e+07u w=1.72e+07u
X5816 adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5817 adc_array_wafflecap_8_8_0[12|8]/adc_array_circuit_150n_0/vint2 row_n[8] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5818 adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5819 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vint1 row_n[20] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5820 adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5821 adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5822 adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5823 VDD VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5824 VSS col_n[1] adc_array_wafflecap_8_8_0[1|25]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5825 adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5826 adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5827 adc_array_wafflecap_8_8_0[7|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5828 VSS col_n[4] adc_array_wafflecap_8_8_0[4|3]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5829 adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5830 adc_array_wafflecap_8_8_0[14|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5831 adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|4]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5832 VSS col_n[7] adc_array_wafflecap_8_8_0[7|15]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5833 VSS sample_n adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5834 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5835 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5836 adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vdrv col_n[10] adc_array_wafflecap_8_8_0[10|8]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5837 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5838 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vint2 colon_n[10] adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5839 adc_array_wafflecap_8_8_0[8|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5840 adc_array_wafflecap_8_8_0[7|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5841 adc_array_wafflecap_8_8_0[3|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5842 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5843 adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5844 vcom adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5845 adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5846 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5847 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5848 adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5849 adc_array_wafflecap_8_8_0[3|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5850 adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|25]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5851 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5852 adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5853 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vint1 row_n[3] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5854 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5855 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5856 VSS col_n[14] adc_array_wafflecap_8_8_0[14|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5857 VSS col_n[6] adc_array_wafflecap_8_8_0[6|7]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5858 VSS col_n[2] adc_array_wafflecap_8_8_0[2|8]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5859 VSS col_n[13] adc_array_wafflecap_8_8_0[13|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5860 adc_array_wafflecap_8_8_0[15|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5861 adc_array_wafflecap_8_8_0[6|9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5862 adc_array_wafflecap_8_8_0[2|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5863 adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5864 adc_array_wafflecap_8_Dummy_5[14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5865 adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5866 adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5867 VDD VDD adc_array_wafflecap_8_Dummy_4[23]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5868 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5869 adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n sample VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5870 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|26]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5871 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5872 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5873 adc_array_wafflecap_8_8_0[13|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5874 adc_array_wafflecap_8_8_0[12|23]/adc_array_circuit_150n_0/vint1 row_n[23] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5875 VSS col_n[10] adc_array_wafflecap_8_8_0[10|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5876 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5877 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vint1 row_n[8] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5878 VSS col_n[10] adc_array_wafflecap_8_8_0[10|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5879 adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|29]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5880 VSS col_n[11] adc_array_wafflecap_8_8_0[11|6]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5881 adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=1.386e+11p pd=1.5e+06u as=0p ps=0u w=420000u l=150000u
X5882 adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5883 adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[12|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5884 adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vdrv col_n[11] adc_array_wafflecap_8_8_0[11|22]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5885 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|7]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5886 adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5887 vcom VSS adc_array_wafflecap_8_Dummy_0[7]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5888 adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5889 VSS col_n[3] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5890 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint2 colon_n[7] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5891 adc_array_wafflecap_8_8_0[0|2]/adc_array_circuit_150n_0/vint2 row_n[2] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5892 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5893 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5894 VDD colon_n[13] adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5895 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5896 adc_array_wafflecap_8_8_0[13|16]/adc_array_circuit_150n_0/vint2 row_n[16] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5897 adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[11|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5898 adc_array_wafflecap_8_8_0[2|19]/adc_array_circuit_150n_0/vint2 row_n[19] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5899 adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/vint1 row_n[6] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5900 adc_array_wafflecap_8_8_0[15|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5901 adc_array_wafflecap_8_8_0[15|15]/adc_array_circuit_150n_0/vint1 row_n[15] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5902 adc_array_wafflecap_8_8_0[8|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5903 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint2 row_n[9] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5904 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5905 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint2 colon_n[6] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5906 VDD colon_n[5] adc_array_wafflecap_8_8_0[5|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5907 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5908 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5909 adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5910 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5911 adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5912 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5913 adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5914 adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5915 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|2]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5916 adc_array_wafflecap_8_8_0[13|26]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5917 adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5918 adc_array_wafflecap_8_8_0[11|18]/adc_array_circuit_150n_0/vint2 row_n[18] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5919 adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|23]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5920 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5921 VDD colon_n[4] adc_array_wafflecap_8_8_0[4|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5922 adc_array_wafflecap_8_8_0[4|23]/adc_array_circuit_150n_0/vint2 row_n[23] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5923 adc_array_wafflecap_8_Dummy_3[5]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5924 adc_array_wafflecap_8_8_0[0|24]/adc_array_circuit_150n_0/vint2 row_n[24] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5925 vcom adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5926 adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vdrv col_n[8] adc_array_wafflecap_8_8_0[8|9]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5927 adc_array_wafflecap_8_8_0[7|1]/adc_array_circuit_150n_0/vint2 row_n[1] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5928 adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vint2 colon_n[1] adc_array_wafflecap_8_8_0[1|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5929 adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5930 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|9]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5931 adc_array_wafflecap_8_8_0[9|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5932 adc_array_wafflecap_8_8_0[9|13]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5933 adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5934 adc_array_wafflecap_8_8_0[13|17]/adc_array_circuit_150n_0/vint1 row_n[17] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5935 VDD colon_n[11] adc_array_wafflecap_8_8_0[11|21]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5936 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5937 adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vdrv col_n[7] adc_array_wafflecap_8_8_0[7|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5938 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5939 adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vdrv col_n[9] adc_array_wafflecap_8_8_0[9|18]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5940 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vint2 colon_n[9] adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5941 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|8]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5942 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5943 VSS col_n[0] adc_array_wafflecap_8_8_0[0|9]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5944 adc_array_wafflecap_8_8_0[15|30]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5945 adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[13|6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5946 vcom adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5947 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.64e+11p ps=2.26e+06u w=800000u l=150000u
X5948 adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vdrv col_n[2] adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5949 adc_array_wafflecap_8_8_0[14|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5950 vcom adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|3]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5951 adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5952 VDD colon_n[3] adc_array_wafflecap_8_8_0[3|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5953 vcom adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5954 VSS VSS adc_array_wafflecap_8_Dummy_3[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5955 adc_array_wafflecap_8_8_0[2|28]/adc_array_circuit_150n_0/vint2 row_n[28] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5956 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5957 adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vdrv col_n[6] adc_array_wafflecap_8_8_0[6|14]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5958 adc_array_wafflecap_8_8_0[6|27]/adc_array_circuit_150n_0/vint2 row_n[27] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5959 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vint2 VDD adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5960 adc_array_wafflecap_8_8_0[5|6]/adc_array_circuit_150n_0/vint2 row_n[6] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5961 adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|11]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5962 adc_array_wafflecap_8_Dummy_4[20]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5963 VSS col_n[12] adc_array_wafflecap_8_8_0[12|14]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5964 adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vint2 colon_n[2] adc_array_wafflecap_8_8_0[2|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5965 adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5966 adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|15]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5967 VSS col_n[12] adc_array_wafflecap_8_8_0[12|4]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5968 adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[9|27]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5969 VSS col_n[8] adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5970 adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5971 adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5972 adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|27]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5973 adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5974 adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|28]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5975 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|13]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5976 adc_array_wafflecap_8_8_0[11|10]/adc_array_circuit_150n_0/vint1 row_n[10] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5977 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vint2 colon_n[11] adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5978 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5979 VDD colon_n[14] adc_array_wafflecap_8_8_0[14|3]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5980 adc_array_wafflecap_8_8_0[12|18]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5981 adc_array_wafflecap_8_8_0[11|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5982 adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/vint1 row_n[4] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5983 adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/vint1 row_n[14] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5984 VDD colon_n[0] adc_array_wafflecap_8_8_0[0|15]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5985 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5986 vcom adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[13|18]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5987 adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[8|21]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5988 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5989 adc_array_wafflecap_8_8_0[3|18]/adc_array_circuit_150n_0/vint1 row_n[18] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5990 adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|1]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5991 adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5992 adc_array_wafflecap_8_8_0[8|19]/adc_array_circuit_150n_0/vint1 row_n[19] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5993 adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[7|12]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5994 adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[3|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[3|13]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5995 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|29]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5996 adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vdrv col_n[3] adc_array_wafflecap_8_8_0[3|16]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5997 adc_array_wafflecap_8_Dummy_5[0]/adc_array_circuit_150n_0/vint2 VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5998 adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X5999 VDD colon_n[9] adc_array_wafflecap_8_8_0[9|17]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6000 adc_array_wafflecap_8_8_0[9|21]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6001 adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[1|20]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6002 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vint2 colon_n[14] adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6003 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|16]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6004 adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[7|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6005 adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|12]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6006 adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vint2 colon_n[13] adc_array_wafflecap_8_8_0[13|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6007 vcom adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|6]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6008 adc_array_wafflecap_8_Dummy_0[1]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6009 vcom VSS adc_array_wafflecap_8_Dummy_4[30]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6010 adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vdrv col_n[15] adc_array_wafflecap_8_8_0[15|2]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6011 VSS col_n[6] adc_array_wafflecap_8_8_0[6|0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6012 adc_array_wafflecap_8_Dummy_4[25]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6013 VSS col_n[5] adc_array_wafflecap_8_8_0[5|13]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6014 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6015 VSS col_n[10] adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6016 adc_array_wafflecap_8_8_0[6|24]/adc_array_circuit_150n_0/vint1 row_n[24] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6017 adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6018 VDD colon_n[12] adc_array_wafflecap_8_8_0[12|19]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6019 adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[15|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6020 adc_array_wafflecap_8_8_0[13|28]/adc_array_circuit_150n_0/vint1 row_n[28] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6021 VDD colon_n[11] adc_array_wafflecap_8_Dummy_5[11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6022 adc_array_wafflecap_8_8_0[1|22]/adc_array_circuit_150n_0/vint1 row_n[22] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6023 adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[6|2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6024 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|29]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6025 VDD colon_n[1] adc_array_wafflecap_8_Dummy_5[1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6026 adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[2|3]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6027 adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[5|15]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6028 adc_array_wafflecap_8_8_0[4|0]/adc_array_circuit_150n_0/vint1 row_n[0] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6029 adc_array_wafflecap_8_8_0[1|17]/adc_array_circuit_150n_0/vint2 row_n[17] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6030 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6031 adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|10]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6032 adc_array_wafflecap_8_Dummy_2[5]/adc_array_circuit_150n_0/cbot VDD vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6033 VSS col_n[1] adc_array_wafflecap_8_8_0[1|27]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6034 adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[9|0]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6035 adc_array_wafflecap_8_8_0[7|31]/adc_array_circuit_150n_0/vint2 row_n[31] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6036 VSS col_n[4] adc_array_wafflecap_8_8_0[4|5]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6037 VSS VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6038 adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|19]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6039 adc_array_wafflecap_8_Dummy_4[31]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6040 VSS col_n[13] adc_array_wafflecap_8_8_0[13|2]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6041 VSS col_n[13] adc_array_wafflecap_8_8_0[13|12]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6042 adc_array_wafflecap_8_8_0[7|7]/adc_array_circuit_150n_0/vint1 row_n[7] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6043 adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[14]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6044 adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[10|25]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6045 adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/vdrv VSS adc_array_wafflecap_8_Dummy_4[4]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6046 adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vdrv col_n[12] adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6047 adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample sample_n VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6048 adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|26]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6049 adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vdrv col_n[5] adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6050 adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[4|7]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6051 adc_array_wafflecap_8_8_0[3|26]/adc_array_circuit_150n_0/vint1 row_n[26] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6052 adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[0|8]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6053 adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[12|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[12|16]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6054 adc_array_wafflecap_8_8_0[2|5]/adc_array_circuit_150n_0/vint1 row_n[5] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6055 VSS sample adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample_n VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6056 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6057 adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[15|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[15|7]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6058 VDD colon_n[15] adc_array_wafflecap_8_8_0[15|11]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6059 VSS VSS adc_array_wafflecap_8_Dummy_2[0]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6060 adc_array_wafflecap_8_8_0[6|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6061 adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6062 VSS col_n[9] adc_array_wafflecap_8_8_0[9|23]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6063 VDD VSS adc_array_wafflecap_8_Dummy_2[6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6064 adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vint2 colon_n[5] adc_array_wafflecap_8_8_0[5|23]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6065 adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vint2 colon_n[8] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6066 adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|28]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6067 adc_array_wafflecap_8_8_0[10|19]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6068 adc_array_wafflecap_8_Dummy_5[9]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[9|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6069 vcom VSS adc_array_wafflecap_8_Dummy_4[28]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6070 adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6071 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|14]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6072 vcom adc_array_wafflecap_8_8_0[10|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[10|4]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6073 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[4|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6074 adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vint2 colon_n[4] adc_array_wafflecap_8_8_0[4|12]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6075 adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6076 adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[1|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6077 adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[14|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[14|19]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6078 vcom adc_array_wafflecap_8_8_0[11|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[11|8]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6079 VDD colon_n[8] adc_array_wafflecap_8_8_0[8|1]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6080 VDD colon_n[7] adc_array_wafflecap_8_8_0[7|14]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6081 vcom adc_array_wafflecap_8_8_0[0|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[0|19]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6082 adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vint2 colon_n[3] adc_array_wafflecap_8_8_0[3|28]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6083 adc_array_wafflecap_8_8_0[6|20]/adc_array_circuit_150n_0/vint2 row_n[20] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6084 adc_array_wafflecap_8_8_0[2|21]/adc_array_circuit_150n_0/vint2 row_n[21] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6085 VDD colon_n[2] adc_array_wafflecap_8_8_0[2|12]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6086 adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|10]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6087 VSS col_n[6] adc_array_wafflecap_8_8_0[6|30]/adc_array_circuit_150n_0/vint2 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6088 adc_array_wafflecap_8_8_0[15|29]/adc_array_circuit_150n_0/vint2 row_n[29] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6089 adc_array_wafflecap_8_8_0[13|11]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6090 adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vint2 colon_n[12] adc_array_wafflecap_8_8_0[12|0]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6091 adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/vdrv adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|17]/adc_array_circuit_150n_0/cbot VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6092 adc_array_wafflecap_8_8_0[8|11]/adc_array_circuit_150n_0/vint2 row_n[11] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6093 adc_array_wafflecap_8_8_0[13|1]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[13|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6094 adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vdrv col_n[13] adc_array_wafflecap_8_8_0[13|25]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6095 adc_array_wafflecap_8_8_0[8|27]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample_n vcom VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6096 adc_array_wafflecap_8_8_0[11|29]/adc_array_circuit_150n_0/vint1 row_n[29] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6097 VDD colon_n[6] adc_array_wafflecap_8_8_0[6|6]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6098 adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vint2 VSS adc_array_wafflecap_8_Dummy_1[2]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6099 vcom adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[6|22]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6100 vcom adc_array_wafflecap_8_8_0[2|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[2|23]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6101 adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/cbot adc_array_wafflecap_8_8_0[6|31]/adc_array_circuit_150n_0/sample_n adc_array_wafflecap_8_Dummy_5[6]/adc_array_circuit_150n_0/vdrv VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6102 vcom adc_array_wafflecap_8_8_0[5|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[5|1]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6103 adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vdrv col_n[4] adc_array_wafflecap_8_8_0[4|20]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6104 adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vdrv col_n[0] adc_array_wafflecap_8_8_0[0|21]/adc_array_circuit_150n_0/vint1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6105 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|10]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6106 vcom adc_array_wafflecap_8_8_0[8|31]/adc_array_circuit_150n_0/sample adc_array_wafflecap_8_8_0[8|13]/adc_array_circuit_150n_0/cbot VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6107 adc_array_wafflecap_8_8_0[4|30]/adc_array_circuit_150n_0/vint1 row_n[30] VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6108 VDD colon_n[1] adc_array_wafflecap_8_8_0[1|4]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6109 VDD colon_n[10] adc_array_wafflecap_8_8_0[10|0]/adc_array_circuit_150n_0/vdrv VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=800000u l=150000u
X6110 adc_array_wafflecap_8_8_0[4|25]/adc_array_circuit_150n_0/vint2 row_n[25] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6111 adc_array_wafflecap_8_8_0[0|26]/adc_array_circuit_150n_0/vint2 row_n[26] VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

