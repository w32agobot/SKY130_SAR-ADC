magic
tech sky130A
timestamp 1661512818
<< poly >>
rect 0 98 64 114
<< locali >>
rect 44 313 467 330
rect 27 270 57 287
rect 216 119 240 122
rect 216 102 220 119
rect 237 102 240 119
rect 216 98 240 102
rect 464 98 481 118
rect 41 0 367 17
<< viali >>
rect 280 276 297 293
rect 220 102 237 119
<< metal1 >>
rect -3 296 58 299
rect -3 293 303 296
rect -3 282 280 293
rect 272 276 280 282
rect 297 276 303 293
rect 272 273 303 276
rect 42 131 195 149
rect 177 75 195 131
rect 222 131 264 149
rect 324 132 483 150
rect 222 125 240 131
rect 216 119 240 125
rect 216 102 220 119
rect 237 102 240 119
rect 216 96 240 102
rect 177 57 269 75
use NOR  NOR_0 ../NOR
timestamp 1661511935
transform 1 0 4 0 1 118
box -4 -118 253 230
use NOR  NOR_1
timestamp 1661511935
transform 1 0 252 0 1 118
box -4 -118 253 230
<< labels >>
rlabel poly 0 98 0 114 7 R
port 1 w
rlabel metal1 -3 283 -3 299 7 S
port 7 w
rlabel locali 41 0 41 17 7 VSS
port 5 w
rlabel locali 44 313 44 330 7 VDD
port 4 w
rlabel locali 481 98 481 118 3 QN
port 2 e
rlabel metal1 483 132 483 150 3 Q
port 6 e
<< end >>
