magic
tech sky130A
magscale 1 2
timestamp 1665671751
<< nwell >>
rect 141 880 859 1004
rect 0 506 1004 880
rect 141 499 859 506
<< nmos >>
rect 239 51 279 431
rect 337 51 377 431
rect 435 51 475 431
rect 533 51 573 431
rect 631 51 671 431
rect 729 51 769 431
<< pmos >>
rect 235 588 275 968
rect 333 588 373 968
rect 431 588 471 968
rect 529 588 569 968
rect 627 588 667 968
rect 725 588 765 968
<< ndiff >>
rect 181 419 239 431
rect 181 63 193 419
rect 227 63 239 419
rect 181 51 239 63
rect 279 419 337 431
rect 279 63 291 419
rect 325 63 337 419
rect 279 51 337 63
rect 377 419 435 431
rect 377 63 389 419
rect 423 63 435 419
rect 377 51 435 63
rect 475 419 533 431
rect 475 63 487 419
rect 521 63 533 419
rect 475 51 533 63
rect 573 419 631 431
rect 573 63 585 419
rect 619 63 631 419
rect 573 51 631 63
rect 671 419 729 431
rect 671 63 683 419
rect 717 63 729 419
rect 671 51 729 63
rect 769 419 827 431
rect 769 63 781 419
rect 815 63 827 419
rect 769 51 827 63
<< pdiff >>
rect 177 956 235 968
rect 177 600 189 956
rect 223 600 235 956
rect 177 588 235 600
rect 275 956 333 968
rect 275 600 287 956
rect 321 600 333 956
rect 275 588 333 600
rect 373 956 431 968
rect 373 600 385 956
rect 419 600 431 956
rect 373 588 431 600
rect 471 956 529 968
rect 471 607 483 956
rect 517 607 529 956
rect 471 588 529 607
rect 569 956 627 968
rect 569 600 581 956
rect 615 600 627 956
rect 569 588 627 600
rect 667 956 725 968
rect 667 600 679 956
rect 713 600 725 956
rect 667 588 725 600
rect 765 956 823 968
rect 765 600 777 956
rect 811 600 823 956
rect 765 588 823 600
<< ndiffc >>
rect 193 63 227 419
rect 291 63 325 419
rect 389 63 423 419
rect 487 63 521 419
rect 585 63 619 419
rect 683 63 717 419
rect 781 63 815 419
<< pdiffc >>
rect 189 600 223 956
rect 287 600 321 956
rect 385 600 419 956
rect 483 607 517 956
rect 581 600 615 956
rect 679 600 713 956
rect 777 600 811 956
<< poly >>
rect 235 968 275 994
rect 333 968 373 994
rect 431 968 471 994
rect 529 968 569 994
rect 627 968 667 994
rect 725 968 765 994
rect 235 572 275 588
rect 333 572 373 588
rect 235 542 373 572
rect 431 573 471 588
rect 529 573 569 588
rect 627 573 667 588
rect 725 573 765 588
rect 431 543 765 573
rect 239 476 373 542
rect 631 476 765 543
rect 239 446 573 476
rect 239 431 279 446
rect 337 431 377 446
rect 435 431 475 446
rect 533 431 573 446
rect 631 446 769 476
rect 631 431 671 446
rect 729 431 769 446
rect 239 4 279 51
rect 337 4 377 51
rect 435 4 475 51
rect 533 4 573 51
rect 631 4 671 51
rect 729 4 769 51
<< locali >>
rect 34 924 148 1004
rect 34 888 46 924
rect 136 888 148 924
rect 34 706 148 888
rect 34 670 46 706
rect 136 670 148 706
rect 34 610 148 670
rect 34 574 46 610
rect 136 574 148 610
rect 34 266 148 574
rect 34 232 114 266
rect 34 102 148 232
rect 34 66 46 102
rect 136 66 148 102
rect 34 0 148 66
rect 182 956 229 972
rect 182 600 189 956
rect 223 600 229 956
rect 182 419 229 600
rect 277 956 331 972
rect 277 941 287 956
rect 277 897 286 941
rect 277 600 287 897
rect 321 600 331 956
rect 277 572 331 600
rect 374 956 430 972
rect 374 600 385 956
rect 419 600 430 956
rect 374 584 430 600
rect 483 956 517 972
rect 483 591 517 607
rect 581 956 615 972
rect 679 956 713 972
rect 615 630 638 707
rect 581 584 615 600
rect 679 584 713 600
rect 777 956 811 972
rect 777 584 811 600
rect 854 924 970 1004
rect 854 888 866 924
rect 958 888 970 924
rect 854 706 970 888
rect 854 670 866 706
rect 958 670 970 706
rect 854 610 970 670
rect 854 574 866 610
rect 958 574 970 610
rect 182 63 193 419
rect 227 63 229 419
rect 182 47 229 63
rect 280 419 335 435
rect 280 56 291 419
rect 325 56 335 419
rect 280 47 335 56
rect 378 419 434 435
rect 378 63 389 419
rect 423 63 434 419
rect 378 47 434 63
rect 487 419 521 437
rect 487 47 521 56
rect 585 419 619 437
rect 683 419 717 435
rect 619 283 636 345
rect 781 419 815 435
rect 585 47 619 63
rect 683 47 717 63
rect 781 47 815 63
rect 854 340 970 574
rect 854 282 866 340
rect 958 282 970 340
rect 854 102 970 282
rect 854 66 866 102
rect 958 66 970 102
rect 854 0 970 66
<< viali >>
rect 46 888 136 924
rect 46 670 136 706
rect 46 574 136 610
rect 114 232 148 266
rect 46 66 136 102
rect 189 897 223 945
rect 286 897 287 941
rect 287 897 321 941
rect 287 663 321 705
rect 385 893 419 941
rect 483 663 517 705
rect 581 894 615 942
rect 581 645 615 686
rect 777 896 811 944
rect 866 888 958 924
rect 866 670 958 706
rect 866 574 958 610
rect 193 300 227 337
rect 291 63 325 98
rect 291 56 325 63
rect 389 300 423 337
rect 487 63 521 98
rect 487 56 521 63
rect 585 283 619 339
rect 683 300 717 338
rect 780 300 781 338
rect 781 300 814 338
rect 866 282 958 340
rect 866 66 958 102
<< metal1 >>
rect 34 924 148 1004
rect 34 888 46 924
rect 136 888 148 924
rect 34 882 148 888
rect 177 945 817 956
rect 177 897 189 945
rect 223 944 817 945
rect 223 942 777 944
rect 223 941 581 942
rect 223 897 286 941
rect 321 897 385 941
rect 177 893 385 897
rect 419 894 581 941
rect 615 896 777 942
rect 811 896 817 944
rect 615 894 817 896
rect 419 893 817 894
rect 177 882 817 893
rect 854 924 970 1004
rect 854 888 866 924
rect 958 888 970 924
rect 854 882 970 888
rect 0 798 1004 854
rect 0 740 1004 770
rect 34 706 148 712
rect 34 670 46 706
rect 136 670 148 706
rect 34 610 148 670
rect 266 711 530 712
rect 266 659 272 711
rect 324 705 530 711
rect 324 663 483 705
rect 517 663 530 705
rect 854 706 970 712
rect 324 659 530 663
rect 266 656 530 659
rect 569 691 628 704
rect 569 639 571 691
rect 623 639 628 691
rect 569 628 628 639
rect 854 670 866 706
rect 958 670 970 706
rect 34 574 46 610
rect 136 574 148 610
rect 34 568 148 574
rect 854 610 970 670
rect 854 574 866 610
rect 958 574 970 610
rect 854 568 970 574
rect 0 512 1004 540
rect 0 430 1004 458
rect 0 374 1004 402
rect 181 339 826 345
rect 181 337 574 339
rect 181 300 193 337
rect 227 300 389 337
rect 423 300 574 337
rect 181 294 574 300
rect 568 283 574 294
rect 630 338 826 339
rect 630 300 683 338
rect 717 300 780 338
rect 814 300 826 338
rect 630 294 826 300
rect 854 340 970 346
rect 630 283 639 294
rect 108 266 154 278
rect 568 277 639 283
rect 854 282 866 340
rect 958 282 970 340
rect 854 276 970 282
rect 108 248 114 266
rect 0 232 114 248
rect 148 248 154 266
rect 148 232 1004 248
rect 0 220 1004 232
rect 0 136 1004 192
rect 34 102 148 108
rect 34 66 46 102
rect 136 66 148 102
rect 34 0 148 66
rect 266 56 272 108
rect 324 104 330 108
rect 324 98 533 104
rect 325 56 487 98
rect 521 56 533 98
rect 266 47 533 56
rect 854 102 970 108
rect 854 66 866 102
rect 958 66 970 102
rect 285 0 325 47
rect 854 0 970 66
<< via1 >>
rect 272 705 324 711
rect 272 663 287 705
rect 287 663 321 705
rect 321 663 324 705
rect 272 659 324 663
rect 571 686 623 691
rect 571 645 581 686
rect 581 645 615 686
rect 615 645 623 686
rect 571 639 623 645
rect 574 283 585 339
rect 585 283 619 339
rect 619 283 630 339
rect 272 98 324 108
rect 272 56 291 98
rect 291 56 324 98
<< metal2 >>
rect 32 962 972 972
rect 32 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 972 962
rect 32 866 972 906
rect 32 810 42 866
rect 98 810 330 866
rect 386 810 618 866
rect 674 810 906 866
rect 962 810 972 866
rect 32 770 972 810
rect 32 714 42 770
rect 98 754 906 770
rect 98 714 244 754
rect 352 734 906 754
rect 32 674 244 714
rect 32 618 42 674
rect 98 618 138 674
rect 194 618 244 674
rect 32 578 244 618
rect 32 522 42 578
rect 98 522 244 578
rect 32 482 244 522
rect 32 426 42 482
rect 98 426 244 482
rect 32 386 244 426
rect 32 330 42 386
rect 98 330 138 386
rect 194 330 244 386
rect 32 290 244 330
rect 32 234 42 290
rect 98 234 244 290
rect 32 194 244 234
rect 32 138 42 194
rect 98 138 244 194
rect 32 98 244 138
rect 32 42 42 98
rect 98 42 138 98
rect 194 42 244 98
rect 272 711 324 717
rect 272 108 324 659
rect 272 50 324 56
rect 352 597 537 734
rect 659 714 906 734
rect 962 714 972 770
rect 566 694 629 705
rect 566 638 569 694
rect 625 638 629 694
rect 566 628 629 638
rect 659 674 972 714
rect 659 618 810 674
rect 866 618 906 674
rect 962 618 972 674
rect 659 597 972 618
rect 352 578 972 597
rect 352 522 906 578
rect 962 522 972 578
rect 352 482 972 522
rect 352 426 906 482
rect 962 426 972 482
rect 352 386 972 426
rect 352 379 810 386
rect 352 242 540 379
rect 568 339 639 348
rect 568 283 574 339
rect 630 283 639 339
rect 568 273 639 283
rect 667 330 810 379
rect 866 330 906 386
rect 962 330 972 386
rect 667 290 972 330
rect 667 242 906 290
rect 352 234 906 242
rect 962 234 972 290
rect 352 194 972 234
rect 352 138 906 194
rect 962 138 972 194
rect 352 98 972 138
rect 352 49 714 98
rect 32 32 244 42
rect 650 42 714 49
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 972 98
rect 650 32 972 42
<< via2 >>
rect 42 906 98 962
rect 138 906 194 962
rect 234 906 290 962
rect 330 906 386 962
rect 426 906 482 962
rect 522 906 578 962
rect 618 906 674 962
rect 714 906 770 962
rect 810 906 866 962
rect 906 906 962 962
rect 42 810 98 866
rect 330 810 386 866
rect 618 810 674 866
rect 906 810 962 866
rect 42 714 98 770
rect 42 618 98 674
rect 138 618 194 674
rect 42 522 98 578
rect 42 426 98 482
rect 42 330 98 386
rect 138 330 194 386
rect 42 234 98 290
rect 42 138 98 194
rect 42 42 98 98
rect 138 42 194 98
rect 906 714 962 770
rect 569 691 625 694
rect 569 639 571 691
rect 571 639 623 691
rect 623 639 625 691
rect 569 638 625 639
rect 810 618 866 674
rect 906 618 962 674
rect 906 522 962 578
rect 906 426 962 482
rect 574 283 630 339
rect 810 330 866 386
rect 906 330 962 386
rect 906 234 962 290
rect 906 138 962 194
rect 714 42 770 98
rect 810 42 866 98
rect 906 42 962 98
<< metal3 >>
rect 36 962 968 968
rect 36 906 42 962
rect 98 906 138 962
rect 194 906 234 962
rect 290 906 330 962
rect 386 906 426 962
rect 482 906 522 962
rect 578 906 618 962
rect 674 906 714 962
rect 770 906 810 962
rect 866 906 906 962
rect 962 906 968 962
rect 36 900 968 906
rect 36 866 104 900
rect 36 810 42 866
rect 98 810 104 866
rect 324 866 392 900
rect 36 770 104 810
rect 36 714 42 770
rect 98 714 104 770
rect 164 824 264 840
rect 164 756 180 824
rect 248 756 264 824
rect 164 740 264 756
rect 324 810 330 866
rect 386 810 392 866
rect 36 680 104 714
rect 324 680 392 810
rect 612 866 680 900
rect 612 810 618 866
rect 674 810 680 866
rect 900 866 968 900
rect 612 784 680 810
rect 740 824 840 840
rect 740 756 756 824
rect 824 756 840 824
rect 740 740 840 756
rect 900 810 906 866
rect 962 810 968 866
rect 900 770 968 810
rect 36 674 392 680
rect 36 618 42 674
rect 98 618 138 674
rect 194 618 392 674
rect 36 612 392 618
rect 555 699 642 723
rect 555 635 566 699
rect 630 635 642 699
rect 900 714 906 770
rect 962 714 968 770
rect 900 680 968 714
rect 36 578 104 612
rect 555 611 642 635
rect 772 674 968 680
rect 772 618 810 674
rect 866 618 906 674
rect 962 618 968 674
rect 772 612 968 618
rect 36 522 42 578
rect 98 522 104 578
rect 900 578 968 612
rect 36 482 104 522
rect 36 426 42 482
rect 98 426 104 482
rect 164 536 264 552
rect 164 468 180 536
rect 248 468 264 536
rect 164 452 264 468
rect 740 536 840 552
rect 740 468 756 536
rect 824 468 840 536
rect 740 452 840 468
rect 900 522 906 578
rect 962 522 968 578
rect 900 482 968 522
rect 36 392 104 426
rect 900 426 906 482
rect 962 426 968 482
rect 900 392 968 426
rect 36 386 324 392
rect 36 330 42 386
rect 98 330 138 386
rect 194 330 324 386
rect 776 386 968 392
rect 36 324 324 330
rect 558 342 645 366
rect 36 290 104 324
rect 36 234 42 290
rect 98 234 104 290
rect 558 278 570 342
rect 634 278 645 342
rect 776 330 810 386
rect 866 330 906 386
rect 962 330 968 386
rect 776 324 968 330
rect 36 194 104 234
rect 36 138 42 194
rect 98 138 104 194
rect 164 248 264 264
rect 558 254 645 278
rect 900 290 968 324
rect 164 180 180 248
rect 248 180 264 248
rect 164 164 264 180
rect 740 248 840 264
rect 740 180 756 248
rect 824 180 840 248
rect 740 164 840 180
rect 900 234 906 290
rect 962 234 968 290
rect 900 194 968 234
rect 36 104 104 138
rect 900 138 906 194
rect 962 138 968 194
rect 900 104 968 138
rect 36 98 324 104
rect 36 42 42 98
rect 98 42 138 98
rect 194 42 324 98
rect 36 36 324 42
rect 692 98 968 104
rect 692 42 714 98
rect 770 42 810 98
rect 866 42 906 98
rect 962 42 968 98
rect 692 36 968 42
<< via3 >>
rect 180 756 248 824
rect 756 756 824 824
rect 566 694 630 699
rect 566 638 569 694
rect 569 638 625 694
rect 625 638 630 694
rect 566 635 630 638
rect 180 468 248 536
rect 756 468 824 536
rect 570 339 634 342
rect 570 283 574 339
rect 574 283 630 339
rect 630 283 634 339
rect 570 278 634 283
rect 180 180 248 248
rect 756 180 824 248
<< metal4 >>
rect 184 840 244 934
rect 164 824 264 840
rect 164 820 180 824
rect 70 760 180 820
rect 164 756 180 760
rect 248 820 264 824
rect 248 760 360 820
rect 248 756 264 760
rect 164 740 264 756
rect 184 552 244 740
rect 472 701 532 934
rect 760 840 820 934
rect 740 824 840 840
rect 740 820 756 824
rect 646 760 756 820
rect 740 756 756 760
rect 824 820 840 824
rect 824 760 934 820
rect 824 756 840 760
rect 740 740 840 756
rect 472 699 631 701
rect 472 635 566 699
rect 630 635 631 699
rect 472 631 631 635
rect 164 536 264 552
rect 164 532 180 536
rect 70 472 180 532
rect 164 468 180 472
rect 248 468 264 536
rect 164 452 264 468
rect 184 264 244 452
rect 472 344 532 631
rect 760 552 820 740
rect 740 536 840 552
rect 740 468 756 536
rect 824 532 840 536
rect 824 472 934 532
rect 824 468 840 472
rect 740 452 840 468
rect 472 342 635 344
rect 472 278 570 342
rect 634 278 635 342
rect 472 276 635 278
rect 164 248 264 264
rect 164 244 180 248
rect 70 184 180 244
rect 164 180 180 184
rect 248 180 264 248
rect 164 164 264 180
rect 184 70 244 164
rect 472 48 532 276
rect 760 264 820 452
rect 740 248 840 264
rect 740 180 756 248
rect 824 244 840 248
rect 824 184 934 244
rect 824 180 840 184
rect 740 164 840 180
rect 760 70 820 164
<< comment >>
rect 0 972 32 1004
rect 972 972 1004 1004
rect 0 0 32 32
rect 972 0 1004 32
<< labels >>
rlabel metal1 0 740 0 770 7 sample_n
port 2 w
rlabel metal1 0 512 0 540 7 colon_n
port 3 w
rlabel metal1 0 430 0 458 7 col_n
port 4 w
rlabel metal1 0 374 0 402 7 sample
port 5 w
rlabel metal1 0 220 0 248 7 vcom
port 6 w
rlabel metal1 0 136 0 192 7 VSS
port 7 w
rlabel locali 854 0 970 0 5 row_n
port 8 s
rlabel metal1 0 798 0 854 7 VDD
port 13 w
flabel metal1 285 0 325 22 0 FreeSans 64 0 0 0 analog_in
port 16 nsew
<< end >>
