VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_mm_sc_hd_dlyPoly5ns
  CLASS CORE ;
  FOREIGN sky130_mm_sc_hd_dlyPoly5ns ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SITE unithd ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 1.195 2.000 1.365 2.235 ;
        RECT 1.190 1.805 1.365 2.000 ;
        RECT 8.055 1.625 8.225 2.635 ;
        RECT 9.355 1.480 9.525 2.635 ;
        RECT 9.355 1.310 9.935 1.480 ;
        RECT 9.765 0.345 9.935 1.310 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 1.195 1.895 1.365 2.155 ;
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
        RECT 1.165 1.810 1.395 2.480 ;
        RECT 1.190 1.805 1.365 1.810 ;
    END
  END VPWR
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.685800 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.320 0.905 1.405 ;
        RECT 0.105 1.045 0.905 1.320 ;
        RECT 0.105 0.990 0.375 1.045 ;
        RECT 0.565 0.975 0.905 1.045 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.366000 ;
    ANTENNADIFFAREA 0.361800 ;
    PORT
      LAYER li1 ;
        RECT 9.015 1.140 9.185 2.455 ;
        RECT 10.110 1.155 10.445 1.325 ;
        RECT 9.015 1.050 9.450 1.140 ;
        RECT 8.720 0.965 9.450 1.050 ;
        RECT 10.215 0.965 10.445 1.155 ;
        RECT 8.720 0.880 9.185 0.965 ;
        RECT 8.720 0.345 8.890 0.880 ;
    END
  END out
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.250 1.680 5.080 2.300 ;
        RECT 7.210 1.680 7.380 1.755 ;
        RECT 3.250 0.980 7.380 1.680 ;
        RECT 7.710 1.340 7.880 1.565 ;
        RECT 10.205 1.545 10.375 2.455 ;
        RECT 7.710 1.175 7.930 1.340 ;
        RECT 0.335 0.380 0.505 0.715 ;
        RECT 4.865 0.085 7.380 0.980 ;
        RECT 7.760 0.085 7.930 1.175 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 10.205 1.705 10.375 1.945 ;
        RECT 7.710 1.395 7.880 1.565 ;
        RECT 0.335 0.460 0.505 0.635 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 7.650 1.570 7.910 1.600 ;
        RECT 10.175 1.570 10.405 2.010 ;
        RECT 7.650 1.375 10.405 1.570 ;
        RECT 7.650 1.365 7.910 1.375 ;
        RECT 0.305 0.240 0.535 0.700 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 2.070 11.230 2.910 ;
        RECT -0.190 1.235 4.110 2.070 ;
        RECT 7.780 1.235 11.230 2.070 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.110 1.070 7.780 2.070 ;
        RECT 0.005 -0.085 11.035 1.070 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 2.905 1.445 3.075 2.235 ;
        RECT 5.475 1.870 7.035 2.125 ;
        RECT 8.535 1.625 8.705 2.455 ;
        RECT 9.695 1.915 9.895 2.455 ;
        RECT 10.685 1.625 10.885 2.455 ;
        RECT 8.100 1.010 8.455 1.180 ;
        RECT 4.315 0.290 4.485 0.800 ;
        RECT 8.240 0.345 8.410 0.795 ;
        RECT 9.285 0.345 9.455 0.715 ;
        RECT 10.245 0.345 10.415 0.795 ;
      LAYER mcon ;
        RECT 2.905 1.525 3.075 2.085 ;
        RECT 5.680 1.920 5.860 2.090 ;
        RECT 6.170 1.920 6.350 2.090 ;
        RECT 8.535 1.770 8.705 2.225 ;
        RECT 9.725 2.060 9.895 2.255 ;
        RECT 10.685 1.805 10.855 2.215 ;
        RECT 8.155 1.010 8.375 1.180 ;
        RECT 4.315 0.460 4.485 0.640 ;
        RECT 8.240 0.525 8.410 0.715 ;
        RECT 9.285 0.495 9.455 0.665 ;
        RECT 10.245 0.525 10.415 0.695 ;
      LAYER met1 ;
        RECT 2.865 1.680 5.080 2.300 ;
        RECT 8.505 2.150 10.885 2.290 ;
        RECT 5.620 1.890 6.410 2.120 ;
        RECT 5.905 1.680 6.130 1.890 ;
        RECT 8.505 1.710 8.735 2.150 ;
        RECT 9.695 2.000 9.925 2.150 ;
        RECT 10.655 1.745 10.885 2.150 ;
        RECT 2.865 1.115 7.480 1.680 ;
        RECT 8.005 1.115 8.455 1.210 ;
        RECT 2.865 0.980 8.455 1.115 ;
        RECT 4.775 0.920 8.455 0.980 ;
        RECT 4.775 0.710 7.480 0.920 ;
        RECT 4.280 0.465 7.480 0.710 ;
        RECT 8.210 0.605 8.440 0.775 ;
        RECT 9.225 0.605 9.515 0.695 ;
        RECT 10.185 0.605 10.475 0.735 ;
        RECT 8.210 0.565 10.475 0.605 ;
        RECT 8.210 0.465 10.445 0.565 ;
        RECT 4.280 0.390 4.700 0.465 ;
  END
END sky130_mm_sc_hd_dlyPoly5ns
END LIBRARY

