* NGSPICE file created from adc_core_digital.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrtp_2 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__inv_2 A Y VPWR VGND VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_2 VPWR VGND A X B VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_2 VGND VPWR Y A B VNB VPB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 B1 A2 X VGND VPWR VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 B Y A VGND VPWR VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_2 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 VPWR a_82_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_646_47# B2 a_82_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_574_369# a_313_47# a_82_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_574_369# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_82_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B2 a_574_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 X a_82_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_82_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_313_47# A2_N a_313_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_313_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_313_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND A2_N a_313_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_82_21# a_313_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND B1 a_646_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__a21oi_4 B1 A2 A1 Y VGND VPWR VNB VPB
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_2 X A1 A2 B1 A3 VGND VPWR VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_4 B C A D X VPWR VGND VNB VPB
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 B X A C VPWR VGND VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR VNB VPB
X0 a_467_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_467_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_467_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_467_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1083_297# A2 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A3 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21# B1 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_889_297# A2 a_1083_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_639_297# A3 a_889_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A2 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_889_297# A3 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_639_297# A4 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A4 a_467_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_1083_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_79_21# A4 a_639_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_467_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_2 X B1 A1 B2 A2 VGND VPWR C1 VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_2 C A X B D VPWR VGND VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_4 X B2 A1 A2 A3 B1 VGND VPWR VNB VPB
X0 a_27_47# B2 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_277_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_549_297# B2 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_739_297# B2 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_739_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_549_297# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_277_297# A3 a_549_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR B1 a_739_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_47# B1 a_549_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_549_297# A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR a_549_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND a_549_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_549_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_549_297# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_549_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_2 B X A VPWR VGND VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__nand2_2 Y A B VGND VPWR VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__and4_2 X C A B D VGND VPWR VNB VPB
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_2 VPWR VGND B1_N A2 A1 Y VNB VPB
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A X VGND VPWR VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_2 A B C_N X VPWR VGND VNB VPB
X0 a_388_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_176_21# a_27_47# a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_472_297# B a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 X B1 A1 A2 VGND VPWR VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 B1 Y A2 A1 VGND VPWR VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_2 X A2 A1 B1 C1 VGND VPWR VNB VPB
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__o22a_2 A2 X B1 A1 B2 VGND VPWR VNB VPB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_8 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 Q RESET_B D CLK VGND VPWR VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_2 A B X C VGND VPWR VNB VPB
X0 VPWR a_30_53# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_30_53# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_30_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_112_297# C a_30_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_30_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_30_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND C a_30_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_184_297# B a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR A a_184_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_2 B2 A2 X B1 C1 A1 VGND VPWR VNB VPB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_2 C A X B D_N VPWR VGND VNB VPB
X0 a_176_21# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND D_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_555_297# C a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_176_21# a_27_53# a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_387_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_483_297# B a_387_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_27_53# a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR D_N a_27_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_2 B2 B1 Y A1 A2 VGND VPWR VNB VPB
X0 Y B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A1 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y A2 a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_2 B1_N Y A2 A1 VGND VPWR VNB VPB
X0 a_397_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1_N a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y A2 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A1 a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y a_28_297# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_28_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_397_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_229_47# a_28_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y a_28_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_229_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_229_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A1 a_397_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_2 VGND VPWR X C1 B1 A1 A2 A3 VNB VPB
X0 a_79_21# C1 a_635_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_417_47# A2 a_319_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_79_21# A1 a_417_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_319_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_319_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_319_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_635_297# B1 a_319_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 X B2 B1 VPWR VGND VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_2 X B1 A3 A1 A2 VGND VPWR VNB VPB
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 B1 A2 A1 Y VGND VPWR VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N X A2_N B2 B1 VGND VPWR VNB VPB
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_4 A1 B1 C1 B2 X A2 VPWR VGND VNB VPB
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 C Y A B VGND VPWR VNB VPB
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_4 A C B Y VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 Y A B VGND VPWR VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_4 A C Y D B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_4 A2 A1 C1 Y B1 VPWR VGND VNB VPB
X0 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_949_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y C1 a_949_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_781_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_781_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_1301_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y C1 a_781_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_27_297# B1 a_1301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_2 C1 B1 A2 A1 X VPWR VGND VNB VPB
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_2 A Y B C VGND VPWR VNB VPB
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 Y C1 VGND VPWR VNB VPB
X0 a_286_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_286_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A2 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_487_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_286_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A1 a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_487_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_286_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_2 VPWR VGND X B A VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_2 B1_N A1 X A2 VGND VPWR VNB VPB
X0 VGND B1_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_478_47# a_27_93# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_478_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A1 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B1_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_574_297# A2 a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_174_21# a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_2 B1_N A2 X A1 VGND VPWR VNB VPB
X0 VPWR A1 a_485_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_485_297# a_297_93# a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_581_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_21# a_297_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_297_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_485_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_2 X A2 A3 A1 B1 C1 VPWR VGND VNB VPB
X0 X a_91_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_91_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_360_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR B1 a_91_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_360_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_360_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_91_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_91_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_91_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_677_47# B1 a_360_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_460_297# A2 a_360_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_91_21# C1 a_677_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_91_21# A3 a_460_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_2 B1 B2 A3 A2 A1 X VGND VPWR VNB VPB
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_2 B2 X A2 A3 A1 B1 VGND VPWR VNB VPB
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_4 VGND VPWR C1 A1 A2 A3 X B1 VNB VPB
X0 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_861_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1059_47# A2 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_1059_47# A1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A3 a_861_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_109_47# A1 a_1059_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_109_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VPWR A3 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_277_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_109_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_861_47# A2 a_1059_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_4 Q D VPWR SET_B CLK VGND VNB VPB
X0 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_1028_413# a_1598_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X4 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1224_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1296_47# a_1178_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND a_1028_413# a_1598_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_2 VGND VPWR A_N C B_N X D VNB VPB
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_2 D1 A1 B1 C1 X A2 VGND VPWR VNB VPB
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 Y B1 A3 A2 VGND VPWR VNB VPB
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4bb_2 D C B_N A_N Y VGND VPWR VNB VPB
X0 VPWR a_193_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND D a_781_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_193_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_591_47# C a_781_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_781_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_781_47# C a_591_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_193_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y a_193_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_591_47# a_27_47# a_341_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_341_47# a_193_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_341_47# a_27_47# a_591_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_193_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_4 X A B VGND VPWR VNB VPB
X0 a_121_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_35_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_4 Y B A VGND VPWR VNB VPB
X0 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_820_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_902_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y a_38_297# a_902_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_902_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y B a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_820_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_902_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR A a_820_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 Y A VPWR VGND VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 Y A B VGND VPWR VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 Y VGND VPWR VNB VPB
X0 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A2 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1163_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# B1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_803_47# B1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1163_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 Y A2 a_1163_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_445_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_803_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_803_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VGND A1 a_803_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_2 B1 A1 X A2 A4 A3 VGND VPWR VNB VPB
X0 a_381_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A2 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_465_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_381_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A4 a_381_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# A1 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 LO HI VPB VNB VGND VPWR
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__and3b_2 VGND VPWR B X A_N C VNB VPB
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_2 Y C A_N B VGND VPWR VNB VPB
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_4 Y B1 A1 A3 A2 VPWR VGND VNB VPB
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_4 Y A1 B1_N A2 VGND VPWR VNB VPB
X0 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_223_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_658_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_223_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND B1_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_223_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_658_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A2 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y A1 a_658_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y a_27_47# a_223_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_4 A1 X C1 A2 B1 VGND VPWR VNB VPB
X0 VGND A1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_1122_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_950_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_557_47# B1 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_474_47# B1 a_748_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_474_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_79_21# C1 a_557_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_474_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_748_47# C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_474_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_79_21# A2 a_950_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_1122_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_4 X B A VGND VPWR VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_806_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X B a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_806_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_806_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR B a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_806_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_112_47# a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_806_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 VPWR A a_806_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_4 A3 A2 A1 Y B1 VGND VPWR VNB VPB
X0 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A3 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_449_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_31_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_31_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A2 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_27_297# A2 a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A3 a_31_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_31_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_449_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_31_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_2 VPWR VGND X A_N D C B VNB VPB
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_4 Y B1 A2 A1 VPWR VGND VNB VPB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_4 X B1 A3 A2 A1 VGND VPWR VNB VPB
X0 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_2 A B_N X VPWR VGND VNB VPB
X0 VPWR A a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_218_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_300_297# a_27_53# a_218_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_218_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_218_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_218_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_218_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_218_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_2 VPWR VGND X B A_N VNB VPB
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 Y A B C VGND VPWR VNB VPB
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311oi_4 Y B1 A1 A3 C1 A2 VPWR VGND VNB VPB
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_1139_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_109_297# B1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_1139_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y C1 a_1139_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X38 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_4 VGND VPWR C1 B1 X A2 A1 VNB VPB
X0 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_473_297# B1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1123_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_555_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A2 a_1123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_951_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_79_204# A1 a_951_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_79_204# C1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_727_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_2 A3 B1 Y A1 A2 VPWR VGND VNB VPB
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A X VGND VPWR VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR A1 A0 S X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_4 B1 A2 A3 A1 X VGND VPWR VNB VPB
X0 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_277_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_277_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_361_47# A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A3 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X a_277_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_277_47# A1 a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_445_47# A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR a_277_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_277_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_4 C1 A1 A2 B1 B2 X VGND VPWR VNB VPB
X0 a_27_47# B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_47# A2 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_717_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_277_297# B2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# B2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_277_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_277_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47# C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47# B2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_277_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_277_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_109_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_717_297# A2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_109_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_4 A2 A1 X B1 VGND VPWR VNB VPB
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_4 A1 Y A2 B1 B2 VGND VPWR VNB VPB
X0 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_33_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_33_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_797_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B1 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_33_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_797_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y B2 a_797_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 Y B2 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y B1 a_33_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_33_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_4 B A_N Y VGND VPWR VNB VPB
X0 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_2 B A Y D C VGND VPWR VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VPWR VGND VNB VPB
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221oi_2 B2 C1 A2 A1 B1 Y VGND VPWR VNB VPB
X0 Y B1 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_301_297# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_301_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B2 a_383_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A1 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# B2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_735_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_301_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR A2 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_383_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_383_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_735_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_301_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_735_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B1 a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_4 A X B C VPWR VGND VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_109_297# C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_4 D1 C1 B1 A2 A1 Y VGND VPWR VNB VPB
X0 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y D1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_28_297# C1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_1205_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_821_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y A1 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_28_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_455_297# B1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1205_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND A2 a_1205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VPWR A1 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_821_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VPWR A2 a_821_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_455_297# C1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_821_297# B1 a_455_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4b_4 D_N B C A X VGND VPWR VNB VPB
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_215_297# a_109_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR A a_487_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_215_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_487_297# B a_403_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_403_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_215_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_297_297# a_109_93# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_4 A B C_N X VGND VPWR VNB VPB
X0 a_176_21# a_27_47# a_626_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_626_297# B a_542_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_542_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_176_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_176_21# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_176_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_176_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_176_21# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_176_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B a_176_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND C_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211oi_2 A2 C1 B1 Y A1 VPWR VGND VNB VPB
X0 VGND A2 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_37_297# B1 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_485_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_292_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_485_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_37_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A1 a_485_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y C1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_292_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_292_297# B1 a_37_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 B1 A2 C1 Y VGND VPWR VNB VPB
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_4 A_N X C B VGND VPWR VNB VPB
X0 a_98_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_98_199# a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_257_47# B a_152_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_152_47# a_98_199# a_56_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR C a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_98_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_56_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND C a_257_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221ai_2 B1 B2 Y A2 A1 C1 VGND VPWR VNB VPB
X0 Y A2 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_300_47# B2 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_300_47# B1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_734_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_28_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C1 a_28_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_382_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_28_47# B1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_28_47# B2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B2 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_734_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A2 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_382_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_734_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_4 B1_N A1 A2 X VGND VPWR VNB VPB
X0 VPWR B1_N a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_743_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_575_47# a_27_297# a_187_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_743_297# A2 a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_27_297# a_187_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_187_21# A2 a_743_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_187_21# a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_187_21# a_27_297# a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B1_N a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A2 a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A1 a_575_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR a_187_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_575_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_575_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_187_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 X a_187_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND a_187_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_4 X A1 A2 C1 B1 D1 VPWR VGND VNB VPB
X0 VGND A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# A2 a_852_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_852_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_361_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR C1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND A2 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47# D1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_361_47# B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_361_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_277_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_445_47# B1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_681_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_27_47# C1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR D1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A1 a_681_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_27_297# D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4bb_2 A X B D_N C_N VPWR VGND VNB VPB
X0 a_398_413# a_206_93# a_316_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR a_316_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_316_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_316_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_27_410# a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_316_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_316_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_566_297# B a_494_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_206_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_316_413# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_206_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_494_297# a_27_410# a_398_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_316_413# a_206_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VPWR A a_566_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_2 C D Y A B VGND VPWR VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_4 C A_N D X B_N VGND VPWR VNB VPB
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_174_21# a_832_21# a_766_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_832_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_766_47# a_27_47# a_652_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_652_47# C a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_832_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_556_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR a_832_21# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND B_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_2 D1 C1 A2 A1 B1 X VGND VPWR VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt adc_core_digital VGND VPWR clk_dig_in comparator_in config_1_in[0] config_1_in[10]
+ config_1_in[11] config_1_in[12] config_1_in[13] config_1_in[14] config_1_in[15]
+ config_1_in[1] config_1_in[2] config_1_in[3] config_1_in[4] config_1_in[5] config_1_in[6]
+ config_1_in[7] config_1_in[8] config_1_in[9] config_2_in[0] config_2_in[10] config_2_in[11]
+ config_2_in[12] config_2_in[13] config_2_in[14] config_2_in[15] config_2_in[1] config_2_in[2]
+ config_2_in[3] config_2_in[4] config_2_in[5] config_2_in[6] config_2_in[7] config_2_in[8]
+ config_2_in[9] conv_finished_out enable_loop_out nmatrix_bincap_out_n[0] nmatrix_bincap_out_n[1]
+ nmatrix_bincap_out_n[2] nmatrix_c0_out_n nmatrix_col_out_n[0] nmatrix_col_out_n[10]
+ nmatrix_col_out_n[11] nmatrix_col_out_n[12] nmatrix_col_out_n[13] nmatrix_col_out_n[14]
+ nmatrix_col_out_n[15] nmatrix_col_out_n[16] nmatrix_col_out_n[17] nmatrix_col_out_n[18]
+ nmatrix_col_out_n[19] nmatrix_col_out_n[1] nmatrix_col_out_n[20] nmatrix_col_out_n[21]
+ nmatrix_col_out_n[22] nmatrix_col_out_n[23] nmatrix_col_out_n[24] nmatrix_col_out_n[25]
+ nmatrix_col_out_n[26] nmatrix_col_out_n[27] nmatrix_col_out_n[28] nmatrix_col_out_n[29]
+ nmatrix_col_out_n[2] nmatrix_col_out_n[30] nmatrix_col_out_n[31] nmatrix_col_out_n[3]
+ nmatrix_col_out_n[4] nmatrix_col_out_n[5] nmatrix_col_out_n[6] nmatrix_col_out_n[7]
+ nmatrix_col_out_n[8] nmatrix_col_out_n[9] nmatrix_row_out_n[0] nmatrix_row_out_n[10]
+ nmatrix_row_out_n[11] nmatrix_row_out_n[12] nmatrix_row_out_n[13] nmatrix_row_out_n[14]
+ nmatrix_row_out_n[15] nmatrix_row_out_n[1] nmatrix_row_out_n[2] nmatrix_row_out_n[3]
+ nmatrix_row_out_n[4] nmatrix_row_out_n[5] nmatrix_row_out_n[6] nmatrix_row_out_n[7]
+ nmatrix_row_out_n[8] nmatrix_row_out_n[9] nmatrix_rowon_out_n[0] nmatrix_rowon_out_n[10]
+ nmatrix_rowon_out_n[11] nmatrix_rowon_out_n[12] nmatrix_rowon_out_n[13] nmatrix_rowon_out_n[14]
+ nmatrix_rowon_out_n[15] nmatrix_rowon_out_n[1] nmatrix_rowon_out_n[2] nmatrix_rowon_out_n[3]
+ nmatrix_rowon_out_n[4] nmatrix_rowon_out_n[5] nmatrix_rowon_out_n[6] nmatrix_rowon_out_n[7]
+ nmatrix_rowon_out_n[8] nmatrix_rowon_out_n[9] pmatrix_bincap_out_n[0] pmatrix_bincap_out_n[1]
+ pmatrix_bincap_out_n[2] pmatrix_c0_out_n pmatrix_col_out_n[0] pmatrix_col_out_n[10]
+ pmatrix_col_out_n[11] pmatrix_col_out_n[12] pmatrix_col_out_n[13] pmatrix_col_out_n[14]
+ pmatrix_col_out_n[15] pmatrix_col_out_n[16] pmatrix_col_out_n[17] pmatrix_col_out_n[18]
+ pmatrix_col_out_n[19] pmatrix_col_out_n[1] pmatrix_col_out_n[20] pmatrix_col_out_n[21]
+ pmatrix_col_out_n[22] pmatrix_col_out_n[23] pmatrix_col_out_n[24] pmatrix_col_out_n[25]
+ pmatrix_col_out_n[26] pmatrix_col_out_n[27] pmatrix_col_out_n[28] pmatrix_col_out_n[29]
+ pmatrix_col_out_n[2] pmatrix_col_out_n[30] pmatrix_col_out_n[31] pmatrix_col_out_n[3]
+ pmatrix_col_out_n[4] pmatrix_col_out_n[5] pmatrix_col_out_n[6] pmatrix_col_out_n[7]
+ pmatrix_col_out_n[8] pmatrix_col_out_n[9] pmatrix_row_out_n[0] pmatrix_row_out_n[10]
+ pmatrix_row_out_n[11] pmatrix_row_out_n[12] pmatrix_row_out_n[13] pmatrix_row_out_n[14]
+ pmatrix_row_out_n[15] pmatrix_row_out_n[1] pmatrix_row_out_n[2] pmatrix_row_out_n[3]
+ pmatrix_row_out_n[4] pmatrix_row_out_n[5] pmatrix_row_out_n[6] pmatrix_row_out_n[7]
+ pmatrix_row_out_n[8] pmatrix_row_out_n[9] pmatrix_rowon_out_n[0] pmatrix_rowon_out_n[10]
+ pmatrix_rowon_out_n[11] pmatrix_rowon_out_n[12] pmatrix_rowon_out_n[13] pmatrix_rowon_out_n[14]
+ pmatrix_rowon_out_n[15] pmatrix_rowon_out_n[1] pmatrix_rowon_out_n[2] pmatrix_rowon_out_n[3]
+ pmatrix_rowon_out_n[4] pmatrix_rowon_out_n[5] pmatrix_rowon_out_n[6] pmatrix_rowon_out_n[7]
+ pmatrix_rowon_out_n[8] pmatrix_rowon_out_n[9] result_out[0] result_out[10] result_out[11]
+ result_out[12] result_out[13] result_out[14] result_out[15] result_out[1] result_out[2]
+ result_out[3] result_out[4] result_out[5] result_out[6] result_out[7] result_out[8]
+ result_out[9] rst_n sample_matrix_out sample_matrix_out_n sample_switch_out sample_switch_out_n
X_2037_ _2037_/Q fanout170/X _2037_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_2106_ VPWR VGND _2106_/X _2106_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_54_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1270_ _1749_/C _1729_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1606_ VPWR VGND _1606_/A _1897_/A _1626_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_0985_ VGND VPWR _1145_/B _1123_/A _1232_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1537_ _1538_/B _2059_/Q _1538_/C _1537_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1399_ _1729_/A _1406_/C _1399_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1468_ VGND VPWR _1467_/Y _1471_/B _1405_/B _1468_/X _1408_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_2
XFILLER_10_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_269 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1322_ _1321_/Y _1314_/Y _1408_/A _1322_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1253_ _1222_/X _1264_/A _1264_/B _1253_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1184_ _1226_/B _1233_/A _1154_/X _1138_/D _1183_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_0968_ _1997_/Q _1151_/C _1994_/Q _0968_/D _0968_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_15_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1871_ _1869_/X _1513_/S _1870_/X _1871_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1940_ VGND VPWR _2056_/D _1940_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_50_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1305_ _1446_/B _1305_/X _1469_/A _1460_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1236_ _1203_/A _1203_/B _1226_/A _1226_/B _1212_/A _1264_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o41a_4
X_1167_ _1317_/B _1149_/X _1165_/X _1166_/X _1166_/B VGND VPWR _1162_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1098_ _1151_/C _1104_/A _1098_/X _1122_/B _1233_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_20_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1021_ _1148_/A _1020_/X _1262_/B _1262_/C _1238_/C _1019_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_4
X_1785_ VGND VPWR _1988_/D _1785_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1854_ _1906_/A _2026_/D _2006_/D _1854_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1923_ _1923_/B _1923_/X _2022_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1219_ _1219_/A _1219_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_16_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1570_ _1570_/Y _1665_/A _1836_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XANTENNA_5 _1377_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2053_ _2053_/Q fanout167/X _2053_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1004_ VGND VPWR input2/X _0929_/B _1003_/X _1110_/S _1003_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_1768_ _1768_/B _1982_/D _2026_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1906_ _1906_/X _1906_/C _1906_/A _2019_/D _1906_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1837_ VGND VPWR _1929_/S _1836_/X _2009_/D _1837_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1699_ _1840_/C _1751_/B _1861_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_15_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput31 VPWR VGND nmatrix_col_out_n[24] _1461_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput42 VPWR VGND nmatrix_col_out_n[5] _1425_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput75 VPWR VGND nmatrix_rowon_out_n[8] _2082_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput64 VPWR VGND nmatrix_rowon_out_n[11] _2085_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput20 VPWR VGND nmatrix_col_out_n[14] _1443_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput53 VPWR VGND nmatrix_row_out_n[1] _2074_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput86 VPWR VGND pmatrix_col_out_n[15] _1371_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput97 VPWR VGND pmatrix_col_out_n[25] _1398_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1622_ VPWR VGND _2017_/Q _1621_/X _1665_/A _1622_/Y VGND VPWR sky130_fd_sc_hd__a21boi_2
X_1484_ _1644_/B _1869_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
X_1553_ _1553_/A _1612_/B _2061_/Q _1553_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_2036_ _2036_/Q fanout166/X _2036_/D _2039_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_2105_ VGND VPWR _2105_/X _2105_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_270 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0984_ VPWR VGND _1232_/C _2002_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_1536_ _1850_/B _1836_/A _1533_/X _1535_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1605_ _1626_/A _1605_/A _1605_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1467_ _1343_/A _1467_/Y _1409_/B _1469_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1398_ _1398_/X _1460_/B _1408_/B _1396_/Y _1397_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_2019_ _2019_/Q fanout170/X _2019_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_42_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_119 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_99 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1321_ _1409_/B _1405_/B _1343_/A _1321_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1252_ _1222_/X _1264_/B _1242_/A _1252_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_17_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1183_ _1238_/C _1183_/X _1119_/X _1262_/B _1157_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_0967_ VGND VPWR _0968_/D _1995_/Q _1996_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1519_ VPWR VGND _1524_/A _1538_/B _1519_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_15_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_262 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_295 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1870_ _1870_/X _1870_/C _1870_/A _1870_/B _1870_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1235_ _1973_/Q _1235_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1166_ _1166_/B _1166_/X _1166_/A _1166_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1304_ _1460_/B _1350_/B _1390_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_52_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1097_ _1967_/Q _1104_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1999_ _1999_/Q fanout176/X _1999_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_11_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1020_ _1151_/C _1020_/X _1122_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1922_ _2040_/D _1831_/B _2040_/Q _1916_/Y _1921_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1784_ VGND VPWR _1784_/S input7/X _1917_/B _1785_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1853_ _1853_/B _1853_/X _1853_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_6_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1218_ VGND VPWR _1973_/D _1218_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1149_ _1147_/X _1149_/X _1148_/X _1220_/B _1115_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_40_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 _1354_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1003_ _1003_/A _1003_/B _1003_/X _1003_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_2052_ _2052_/Q fanout174/X _2052_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1905_ _2021_/D _1920_/B _1905_/X _1889_/B _1904_/X _2017_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
XFILLER_34_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1767_ VGND VPWR _1768_/B _1982_/Q _1769_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1698_ VPWR VGND _1904_/C _1840_/C _1904_/D VGND VPWR sky130_fd_sc_hd__and2_2
X_1836_ _1836_/C _1836_/A _1836_/X _1836_/B _1839_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
XFILLER_13_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput54 VPWR VGND nmatrix_row_out_n[2] _2075_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput10 VPWR VGND conv_finished_out _2026_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput43 VPWR VGND nmatrix_col_out_n[6] _1426_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput21 VPWR VGND nmatrix_col_out_n[15] _1444_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput32 VPWR VGND nmatrix_col_out_n[25] _1462_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput65 VPWR VGND nmatrix_rowon_out_n[12] _2086_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput76 VPWR VGND nmatrix_rowon_out_n[9] _2083_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput98 VPWR VGND pmatrix_col_out_n[26] _1401_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput87 VPWR VGND pmatrix_col_out_n[16] _1373_/Y VGND VPWR sky130_fd_sc_hd__buf_4
X_1621_ _2064_/Q _1621_/A _1621_/X _2016_/Q _1621_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1552_ VGND VPWR _1552_/S _2014_/Q _1551_/Y _1553_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1483_ _1478_/X _1906_/A _1697_/A _1644_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_2104_ VPWR VGND _2104_/X _2104_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_2035_ _2035_/Q fanout170/X _2035_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_30_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1819_ VPWR VGND _1831_/B _1819_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_26_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_290 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0983_ _2005_/Q _2004_/Q _0988_/B _1232_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1535_ _1535_/Y _2059_/Q _1893_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1604_ _2015_/Q _2062_/Q _1605_/B _2061_/Q _2014_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o22ai_2
X_1397_ _1405_/B _1397_/Y _1423_/A _1706_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21bai_2
X_1466_ VGND VPWR _1466_/X _1408_/A _1460_/Y _1451_/A _1706_/D _1314_/Y VGND VPWR
+ sky130_fd_sc_hd__a311o_2
X_2018_ _2018_/Q fanout171/X _2018_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_18_205 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_96 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1320_ VPWR VGND _1405_/B _1320_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1251_ _1250_/X _1264_/B _1234_/B _1974_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1182_ _1201_/B _1193_/A _1201_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_17_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0966_ _1998_/Q _2001_/Q _1999_/Q _2000_/Q _1151_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1518_ _2010_/Q _2057_/Q _1519_/B _2058_/Q _2011_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1449_ _1449_/X _1366_/X _1451_/B _1451_/A _1446_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_9_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1303_ VPWR VGND _1446_/B _1404_/C VGND VPWR sky130_fd_sc_hd__buf_4
X_1234_ VGND VPWR _1242_/A _1974_/Q _1234_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1165_ _1165_/A _1173_/C _1165_/X _1165_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1096_ _1095_/Y _1094_/Y _1040_/D _1166_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_20_244 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0949_ _2043_/D _2043_/Q _0949_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1998_ _1998_/Q fanout176/X _1998_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_28_322 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1921_ _1920_/X _1928_/B _1921_/X _1919_/X _1858_/A _2017_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1852_ _1853_/B _1850_/Y _2014_/D _1851_/X _1849_/X VGND VPWR _1861_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1783_ VGND VPWR _1987_/D _1783_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1217_ VPWR VGND _2104_/A _1218_/A _1217_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1079_ _1198_/A _1105_/A _1105_/B _1105_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1148_ _1148_/X _1148_/C _1148_/A _1148_/B _1148_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_4_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2051_ _2051_/Q fanout173/X _2051_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1002_ _1001_/X _0997_/X _2066_/Q _1003_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1904_ _1904_/X _1904_/C _1904_/A _1906_/A _1904_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1835_ _1836_/B _1835_/X _1834_/X _1836_/C _1786_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_2
X_1697_ _1904_/D _1697_/C _1697_/A _1697_/B _1697_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1766_ _1864_/A _1769_/B _1981_/Q _1766_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_13_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_144 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput55 VPWR VGND nmatrix_row_out_n[3] _2076_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput44 VPWR VGND nmatrix_col_out_n[7] _1428_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput99 VPWR VGND pmatrix_col_out_n[27] _1402_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput66 VPWR VGND nmatrix_rowon_out_n[13] _2087_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput11 VPWR VGND enable_loop_out _2106_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput77 VPWR VGND pmatrix_bincap_out_n[0] _0993_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput88 VPWR VGND pmatrix_col_out_n[17] _1377_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput33 VPWR VGND nmatrix_col_out_n[26] _1465_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput22 VPWR VGND nmatrix_col_out_n[16] _1445_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_321 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1482_ VPWR VGND _1906_/A _1482_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1620_ _1620_/X _1619_/X _1632_/B _1606_/A _1615_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1551_ _1551_/Y _1870_/A _2014_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_2103_ VGND VPWR _2103_/X _2103_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2034_ _2034_/Q fanout165/X _2034_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1818_ VGND VPWR _2005_/D _1818_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1749_ _1749_/C _1749_/A _1750_/A _1749_/B _1749_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_45_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0982_ VPWR VGND _1232_/B _2003_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1534_ VPWR VGND _1893_/B _1612_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1603_ _1543_/Y _1547_/Y _1602_/X _1538_/C _1606_/A _1545_/X VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a221o_4
X_1465_ _1465_/X _1463_/X _1451_/A _1464_/X _1460_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_2017_ _2017_/Q fanout171/X _2017_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1396_ _1429_/B _1396_/Y _1706_/D _1408_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_53_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_209 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1250_ _1250_/X _1973_/Q _1974_/Q _1234_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1181_ _1262_/C _1181_/C _1181_/B _1201_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_17_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0965_ _1123_/C _0965_/C _1123_/A _1157_/C _0965_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1517_ _2058_/Q _1524_/A _2011_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1448_ VGND VPWR _1448_/X _1448_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1379_ _1379_/X _1386_/B _1381_/B _1749_/A _1404_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_23_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1302_ _1404_/C _1311_/A _1311_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1233_ _1233_/A _1233_/C _1234_/B _1233_/D _1262_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4_4
X_1095_ _0968_/X _0965_/X _1223_/A _1095_/Y _1105_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a211oi_4
X_1164_ _1163_/X _1162_/X _1149_/X _1317_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_20_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1997_ _1997_/Q fanout176/X _1997_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0948_ _0946_/Y _0949_/B _0947_/X _2052_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_18_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1851_ _1929_/S _1829_/B _2008_/D _1917_/B _1851_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1920_ VPWR VGND _2023_/D _1920_/X _1920_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1782_ VGND VPWR _1784_/S input6/X _1929_/S _1783_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1216_ VGND VPWR _1216_/S _1749_/A _1973_/Q _1217_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_1147_ _1148_/A _1148_/B _1147_/X _1148_/D _1148_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1078_ _1105_/A _1211_/A _1105_/B _1105_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_2
XFILLER_43_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2050_ _2050_/Q fanout175/X _2050_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_34_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1001_ _1001_/X _1000_/X _0996_/X _0997_/S input2/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_34_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1765_ _1981_/Q _1882_/A _1981_/D _1764_/X _1751_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1903_ _1917_/B _1877_/A _1829_/B _1903_/Y _1929_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_2
X_1834_ _1834_/X _1882_/A _1839_/A _1836_/C _1869_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1696_ VPWR VGND _1697_/D _1928_/B _1980_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_13_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_189 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput23 VPWR VGND nmatrix_col_out_n[17] _1448_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput12 VPWR VGND nmatrix_bincap_out_n[0] _1007_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput34 VPWR VGND nmatrix_col_out_n[27] _1466_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput45 VPWR VGND nmatrix_col_out_n[8] _1431_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput89 VPWR VGND pmatrix_col_out_n[18] _1380_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput78 VPWR VGND pmatrix_bincap_out_n[1] _1032_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput67 VPWR VGND nmatrix_rowon_out_n[14] _2088_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput56 VPWR VGND nmatrix_row_out_n[4] _2077_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1481_ input8/X input7/X _1482_/A input6/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1550_ _1552_/S _1550_/X _1549_/Y _2014_/Q _1836_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_2033_ _2033_/Q fanout170/X _2033_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_2102_ VGND VPWR _2102_/X _2102_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_47_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1748_ VGND VPWR _2102_/A _1748_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1817_ VGND VPWR _1817_/S _1963_/S _2005_/Q _1818_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1679_ VGND VPWR _1679_/Y _1988_/Q _1984_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_3_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_218 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0981_ VPWR VGND _1144_/A _2000_/Q VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_8_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1602_ _2061_/Q _2014_/Q _1602_/X _2015_/Q _2062_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1533_ _1533_/X _2012_/Q _1531_/Y _1532_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1464_ _1469_/C _1464_/X _1464_/A _1464_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1395_ _1395_/X _1406_/B _1460_/B _1343_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2016_ _2016_/Q fanout171/X _2016_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_41_210 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1180_ _1232_/C _1180_/B _1181_/C _1227_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0964_ _1994_/Q _1995_/Q _1157_/C _1996_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1516_ _2010_/Q _1847_/B _2010_/D _1665_/A _1515_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1447_ _1379_/X _1366_/X _1448_/A _1446_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_2
X_1378_ _1451_/B _1408_/B _1378_/X _1469_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
XFILLER_23_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_243 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1232_ _1232_/C _2005_/Q _1233_/D _1232_/B _2004_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1301_ VPWR VGND _1469_/A _1435_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_52_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1094_ _1156_/A _1233_/A _1094_/Y _1150_/B _1105_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4_4
X_1163_ _1163_/X _1289_/A _1165_/C _1173_/B _1162_/B _1166_/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__o311a_2
XFILLER_20_224 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1996_ _1996_/Q fanout175/X _1996_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0947_ _0947_/B _0947_/X _2051_/Q _0947_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_7_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1781_ VPWR VGND _1929_/S _1987_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1850_ _1917_/B _1850_/Y _1850_/B _1850_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_2
X_1215_ VPWR VGND _1749_/A _1404_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1146_ _0990_/C _1145_/A _1145_/X _1262_/C _1227_/C _1148_/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_1077_ _1150_/B _1123_/A _1105_/C _1156_/A _1077_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1979_ _1979_/Q fanout170/X _1979_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_29_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1000_ _2065_/Q _1000_/X _2052_/Q _0914_/C _2067_/Q _0999_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a32o_2
X_1902_ _2026_/D _2037_/D _1900_/X _2037_/Q _1901_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_19_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1764_ VGND VPWR _1766_/C _1762_/Y _1981_/Q _1764_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1833_ _1923_/B _1987_/Q _1833_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1695_ VPWR VGND _1928_/B _1695_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_25_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_124 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1129_ VGND VPWR _1262_/C _1125_/X _1126_/X _1127_/X _1129_/X _1128_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_4
Xoutput24 VPWR VGND nmatrix_col_out_n[18] _1450_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput57 VPWR VGND nmatrix_row_out_n[5] _2078_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput13 VPWR VGND nmatrix_bincap_out_n[1] _1033_/B VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput46 VPWR VGND nmatrix_col_out_n[9] _1434_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput35 VPWR VGND nmatrix_col_out_n[28] _1468_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput68 VPWR VGND nmatrix_rowon_out_n[1] _2075_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput79 VPWR VGND pmatrix_bincap_out_n[2] _1070_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1480_ _1982_/Q _1986_/Q _1980_/Q _1480_/D _1697_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_2032_ _2032_/Q fanout168/X _2032_/D _2060_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_47_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_2101_ VGND VPWR _2101_/X _2101_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1678_ VPWR VGND _1917_/B _1988_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1747_ _1749_/B _1747_/B _1748_/A _1749_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1816_ VGND VPWR _2004_/D _1816_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0980_ VPWR VGND _1262_/C _0980_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_8_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1601_ VPWR VGND _1893_/A _2016_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1532_ _1532_/A _1538_/B _1532_/X _1538_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1394_ _1394_/B _1406_/B _1729_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1463_ _1463_/X _1423_/A _1706_/D _1446_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2015_ _2015_/Q fanout171/X _2015_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_299 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_123 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0963_ VGND VPWR _0965_/C _1997_/Q _1177_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1515_ _1870_/C _1612_/B _1515_/X _1870_/B _1513_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1446_ _1446_/B _1446_/X _1729_/A _1464_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_55_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1377_ _1375_/Y _1377_/X _1387_/A _1471_/A _1412_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_48_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1231_ _1231_/X _1230_/X _1211_/A _1267_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1162_ _1162_/X _1166_/B _1166_/A _1162_/B _1166_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1300_ VPWR VGND _1409_/B _1706_/D VGND VPWR sky130_fd_sc_hd__buf_6
X_1093_ VPWR VGND _1148_/D _1093_/X _1114_/D VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_9_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1995_ _1995_/Q fanout176/X _1995_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0946_ _0947_/B _0947_/C _2051_/Q _0946_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1429_ _1429_/B _1429_/X _1469_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_11_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1780_ _1780_/B _1986_/D _2026_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_6_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1214_ VPWR VGND _1344_/B _1404_/B _1344_/C VGND VPWR sky130_fd_sc_hd__and2_2
X_1145_ _1150_/B _1145_/A _1145_/X _1145_/B _1145_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1076_ _1122_/B _1122_/C _1077_/D _1122_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1978_ _1978_/Q _1978_/D VPWR fanout165/X _2034_/CLK VGND VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_20_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0929_ _0929_/B _1793_/S _1003_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_29_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_70 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1832_ _2029_/D _1831_/X _1830_/X _2026_/D _1822_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1901_ _1901_/X _1831_/B _1861_/B _2012_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1763_ _1979_/Q _1766_/C _1978_/Q _1980_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1694_ _1988_/Q _1989_/Q _1987_/Q _1695_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_25_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1128_ _2005_/Q _1154_/A _1156_/B _1128_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1059_ VGND VPWR _1991_/Q _1956_/B _1993_/Q _1059_/X _1103_/A VGND VPWR sky130_fd_sc_hd__and4bb_2
XFILLER_40_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput14 VPWR VGND nmatrix_bincap_out_n[2] _1070_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput25 VPWR VGND nmatrix_col_out_n[19] _1453_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput47 VPWR VGND nmatrix_row_out_n[10] _2083_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput36 VPWR VGND nmatrix_col_out_n[29] _1470_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput58 VPWR VGND nmatrix_row_out_n[6] _2079_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput69 VPWR VGND nmatrix_rowon_out_n[2] _2076_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2100_ VGND VPWR _2100_/X _2100_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2031_ _2031_/Q fanout165/X _2031_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1815_ VGND VPWR _1817_/S _2005_/Q _2004_/Q _1816_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1677_ input8/X input6/X input7/X _1861_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_7_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1746_ VGND VPWR _2101_/A _1746_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_5_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_187 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1600_ _1877_/A _2015_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1531_ _1538_/B _1538_/C _1532_/A _1531_/Y _1869_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_2
X_1462_ _1408_/A _1423_/A _1372_/X _1460_/Y _1462_/X _1469_/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_1393_ _1393_/X _1391_/C _1341_/Y _1435_/B _1471_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_2014_ _2014_/Q fanout171/X _2014_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1729_ _1729_/C _1729_/A _1730_/A _1729_/B _1749_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_0962_ VPWR VGND _1177_/B _1998_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_1514_ _2010_/Q _1870_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1445_ _1445_/X _1350_/B _1409_/B _1366_/X _1429_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1376_ _1376_/C _1387_/A _1376_/A _1436_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_14_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1092_ VPWR VGND _1289_/A _1173_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1230_ _1230_/X _1226_/Y _1191_/Y _1229_/X _1201_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1161_ _1160_/X _1166_/C _1967_/Q _1053_/X _1041_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_2
XFILLER_37_326 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1994_ _1994_/Q fanout176/X _1994_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_9_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0945_ _2052_/Q _0947_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1428_ _1428_/X _1419_/Y _1423_/A _1427_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_28_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1359_ _1359_/D _1359_/C _1353_/D _1353_/A _1360_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4bb_2
X_1213_ VGND VPWR _1289_/B _1290_/C _1210_/X _1211_/Y _1344_/C _1219_/A VGND VPWR
+ sky130_fd_sc_hd__a311o_4
X_1144_ _1232_/B _1145_/D _1144_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1075_ _1144_/A _1156_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1977_ _1977_/Q fanout167/X _1977_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0928_ _2047_/Q _0927_/Y _0926_/Y _0929_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_16_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1831_ VPWR VGND _2029_/Q _1831_/X _1831_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1900_ _1899_/X _1895_/X _1889_/B _2020_/D _1900_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1762_ _1882_/A _1762_/Y _1981_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1693_ VPWR VGND _1697_/C _1693_/B _1986_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1127_ _1127_/X _1015_/Y _1014_/Y _1016_/X _1123_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1058_ VGND VPWR _1992_/Q _1160_/A _1057_/Y _1058_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput48 VPWR VGND nmatrix_row_out_n[11] _2084_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput26 VPWR VGND nmatrix_col_out_n[1] _1415_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput15 VPWR VGND nmatrix_col_out_n[0] _1414_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput37 VPWR VGND nmatrix_col_out_n[2] _1417_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput59 VPWR VGND nmatrix_row_out_n[7] _2080_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_12_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2030_ _2030_/Q fanout166/X _2030_/D _2039_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1745_ _1747_/B _1749_/D _1712_/C _1746_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1814_ VGND VPWR _2003_/D _1814_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1676_ VPWR VGND _1977_/D _1956_/D VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_53_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1530_ _2059_/Q _1532_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1461_ _1461_/X _1460_/Y _1423_/A _1429_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1392_ VPWR VGND _1392_/X _1392_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_2013_ _2013_/Q fanout167/X _2013_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1728_ VPWR VGND _2087_/A _1728_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1659_ VGND VPWR _1660_/B _2022_/Q _1659_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_32_279 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0961_ _1123_/C _2001_/Q _2000_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1513_ VGND VPWR _1513_/S _1870_/C _1505_/Y _1513_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1444_ _1412_/B _1337_/X _1435_/B _1444_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1375_ _1366_/X _1451_/B _1343_/A _1375_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_46_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1160_ _1229_/D _1160_/X _1160_/A _1160_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1091_ _1173_/C _1202_/B _1969_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_9_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1993_ _1993_/Q fanout176/X _1993_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0944_ _0944_/B _2051_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1427_ _1429_/B _1427_/X _1446_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1358_ _1359_/D _1404_/C _1386_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1289_ _1290_/D _1289_/A _1289_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_6_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1212_ VPWR VGND _1212_/A _1219_/A _1212_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_37_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1074_ _1105_/A _1968_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_4
X_1143_ _2004_/Q _1227_/C _2005_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_37_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_135 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0927_ _2067_/Q _0927_/Y _0926_/A _0914_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1976_ _1976_/Q fanout175/X _1976_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_3_201 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1761_ _1980_/Q _1882_/A _1980_/D _1760_/X _1751_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1830_ VGND VPWR _1833_/B _1828_/X _2012_/D _1830_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1692_ _1693_/B _1989_/Q _1849_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1126_ _1126_/A _1156_/A _1126_/X _1262_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1057_ _1150_/C _1057_/Y _1150_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1959_ VGND VPWR _1963_/S input3/X _2065_/Q _1960_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput38 VPWR VGND nmatrix_col_out_n[30] _1472_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput49 VPWR VGND nmatrix_row_out_n[12] _2085_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput16 VPWR VGND nmatrix_col_out_n[10] _1437_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput27 VPWR VGND nmatrix_col_out_n[20] _1455_/X VGND VPWR sky130_fd_sc_hd__buf_4
XPHY_100 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1744_ _2100_/A _2081_/A _1744_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_30_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1813_ VGND VPWR _1817_/S _2004_/Q _1232_/B _1814_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1675_ VPWR VGND _1956_/D _1675_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_2089_ VGND VPWR _2089_/X _2089_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1109_ VPWR VGND _1109_/X _1109_/B _1289_/A VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_42_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1391_ _1391_/C _1391_/A _1392_/A _1391_/B _1390_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1460_ _1460_/B _1460_/Y _1749_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_2012_ _2012_/Q fanout168/X _2012_/D _2060_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_50_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1658_ _1659_/B _1671_/B _2020_/Q _2021_/Q _1671_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1727_ _1729_/B _1744_/B _1749_/B _1728_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1589_ _1598_/B _1882_/A _2015_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0960_ VPWR VGND _1123_/A _1999_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_1512_ VPWR VGND _1612_/B _1621_/D VGND VPWR sky130_fd_sc_hd__buf_6
X_1374_ _1435_/B _1344_/C _1344_/B _1451_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1443_ VGND VPWR _1443_/X _1443_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1090_ VPWR VGND _1090_/A _1202_/B _1090_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_9_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1992_ _1992_/Q fanout174/X _1992_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0943_ VGND VPWR _0944_/B _2051_/Q _0947_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1426_ _1426_/X _1343_/A _1423_/A _1370_/X _1424_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1357_ _1386_/B _1399_/A _1390_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_1288_ _1290_/A _1290_/B _1289_/B _1290_/C _1289_/A _1288_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_55_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1142_ _1142_/B _1970_/D _1963_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1211_ _1211_/Y _1211_/A _1211_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_37_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1073_ VGND VPWR _1967_/D _1073_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1975_ _1975_/Q fanout174/X _1975_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0926_ _0926_/Y _0926_/A _0926_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1409_ _1409_/Y _1451_/A _1409_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_16_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1760_ VGND VPWR _1760_/S _1980_/Q _1758_/Y _1760_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1691_ _1478_/X _1915_/B _1982_/Q _1697_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1125_ _1144_/A _1262_/D _1126_/A _1125_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1056_ _1019_/X _1056_/Y _1238_/C _1233_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1889_ _1889_/B _1889_/X _2019_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
Xoutput17 VPWR VGND nmatrix_col_out_n[11] _1438_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput28 VPWR VGND nmatrix_col_out_n[21] _1456_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput39 VPWR VGND nmatrix_col_out_n[31] _1473_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1958_ _1957_/X _2104_/A _2064_/D _1216_/S _1977_/D _1747_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41o_2
XPHY_101 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1743_ _2099_/A _1724_/A _1724_/B _1735_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1812_ VGND VPWR _2002_/D _1812_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1674_ VPWR VGND _1991_/Q _1675_/A _1793_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_2088_ VGND VPWR _2088_/X _2088_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xadc_core_digital_193 nmatrix_c0_out_n adc_core_digital_193/HI VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__conb_1
X_1039_ _1123_/A _1233_/C _1157_/B _1040_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_4
X_1108_ _1109_/B _1108_/A _1108_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_12_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1390_ _1390_/A _1404_/C _1390_/X _1429_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_2011_ _2011_/Q fanout167/X _2011_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1657_ _1784_/S _1656_/X _1655_/X _2021_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1588_ _2062_/Q _1588_/X _1864_/A _1893_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1726_ VGND VPWR _2086_/A _1726_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_193 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1511_ _1511_/B _1847_/B _1836_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1442_ _1364_/X _1366_/X _1443_/A _1436_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_2
X_1373_ _1366_/X _1372_/X _1350_/B _1373_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1709_ VGND VPWR _2081_/A _1710_/A _1733_/A _1744_/B VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_29_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0942_ VPWR VGND _2050_/Q _0947_/C _0942_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1991_ _1991_/Q fanout174/X _1991_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1425_ _1425_/X _1420_/Y _1408_/B _1423_/X _1424_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1356_ _1404_/B _1404_/C _1359_/C _1376_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1287_ _1287_/Y _1289_/A _1289_/B _1290_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3b_2
XFILLER_54_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1141_ VGND VPWR _1259_/B _1399_/A _1154_/A _1142_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_1072_ VPWR VGND _1956_/B _1073_/A _1072_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1210_ _1210_/X _1173_/B _1138_/A _1166_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1974_ _1974_/Q fanout171/X _1974_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_20_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0925_ VGND VPWR _2065_/Q _2046_/Q _0924_/X _0926_/B _2066_/Q VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_1408_ _1408_/Y _1408_/A _1408_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1339_ VPWR VGND _1408_/B _1436_/B VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_3_236 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_302 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1690_ VPWR VGND _1915_/B _1690_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1124_ _2004_/Q _1232_/B _1262_/D _1232_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1055_ _1262_/B _1055_/Y _1233_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1957_ _1957_/X _1956_/X _2064_/Q _1950_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
Xoutput18 VPWR VGND nmatrix_col_out_n[12] _1439_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1888_ _1877_/A _1888_/X _1878_/B _2017_/D _1923_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o2bb2a_2
Xoutput29 VPWR VGND nmatrix_col_out_n[22] _1458_/X VGND VPWR sky130_fd_sc_hd__buf_4
XPHY_102 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_151 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1811_ VGND VPWR _1817_/S _1232_/B _1232_/C _1812_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1673_ _1673_/B _2025_/D _1784_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1742_ _2098_/A _1724_/A _1733_/A _1724_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_26_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xadc_core_digital_194 nmatrix_row_out_n[0] adc_core_digital_194/HI VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
X_2087_ VGND VPWR _2087_/X _2087_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1038_ _1044_/B _1993_/Q _1123_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1107_ _1108_/B _1173_/B _1220_/B _1166_/A _1138_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_4
XFILLER_21_132 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_2010_ _2010_/Q fanout165/X _2010_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1725_ _2081_/A _1744_/B _1735_/C _1726_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1656_ _1656_/C _2021_/Q _1656_/X _1656_/B _2020_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1587_ VPWR VGND _2013_/D _1587_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_49_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1510_ VGND VPWR _1513_/S _1505_/Y _1870_/C _1511_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_1441_ _1441_/Y _1332_/X _1440_/X _1353_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21boi_4
X_1372_ _1404_/C _1372_/X _1729_/A _1457_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1708_ _1749_/B _1733_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
X_1639_ _1784_/S _1637_/Y _1636_/X _2018_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_22_260 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_146 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1990_ _2105_/A _1990_/D VPWR fanout168/X _2060_/CLK VGND VGND VPWR sky130_fd_sc_hd__dfstp_4
X_0941_ _0941_/B _2050_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_13_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1355_ _1376_/C _1435_/A _1355_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1424_ _1424_/X _1278_/A _1731_/A _1412_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_34_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_149 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1286_ _1109_/B _1311_/A _1285_/X _1281_/Y _1283_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o211a_4
X_1140_ _1399_/A _1315_/A _1315_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_8
X_1071_ VGND VPWR _1259_/B _1070_/A _1967_/Q _1072_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_0924_ _2065_/Q _0923_/X _0955_/B _0924_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1973_ _1973_/Q fanout174/X _1973_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1407_ VGND VPWR _1407_/X _1407_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1338_ _1337_/X _1343_/A _1405_/B _1328_/Y _1338_/X _1460_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
XFILLER_24_322 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1269_ _1749_/C _1269_/B _1269_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_51_196 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_215 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_119 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1123_ _1123_/B _1123_/C _1123_/A _1123_/D _1123_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1054_ _1053_/X _1245_/B _1044_/X _1081_/A _1967_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_4
X_1887_ _2013_/D _1858_/A _1928_/B _1887_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1956_ VPWR VGND _1956_/X _1216_/S _1956_/D _1976_/Q _1956_/B VGND VPWR sky130_fd_sc_hd__and4b_2
Xoutput19 VPWR VGND nmatrix_col_out_n[13] _1441_/Y VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_119 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1741_ _2097_/A _1724_/A _1724_/B _1471_/B _1733_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1810_ VGND VPWR _2001_/D _1810_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1672_ VGND VPWR _1673_/B _2025_/Q _1672_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1106_ VPWR VGND _1173_/B _1165_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xadc_core_digital_195 pmatrix_row_out_n[0] adc_core_digital_195/HI VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
X_2086_ VGND VPWR _2086_/X _2086_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1037_ _1963_/S _1992_/Q _1037_/X _1991_/Q _1177_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_42_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1939_ VGND VPWR _1977_/D _1968_/D _2056_/Q _1940_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1724_ _2085_/A _1724_/A _1724_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1655_ _1655_/X _1654_/Y _1671_/C _2020_/Q _1671_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1586_ _1587_/A _1585_/X _1904_/A _1583_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_49_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1371_ _1366_/X _1370_/X _1350_/B _1371_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1440_ _1440_/X _1366_/X _1367_/B _1451_/A _1469_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_23_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1638_ _1784_/S _1836_/A _1869_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_8
X_1707_ VGND VPWR _2074_/A _1707_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1569_ _2011_/Q _1836_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_46_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_176 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0940_ VGND VPWR _0941_/B _2050_/Q _0942_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1354_ VGND VPWR _1354_/X _1354_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1423_ VPWR VGND _1423_/A _1423_/X _1423_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_28_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1285_ _1285_/X _1283_/D _1108_/A _1284_/X _1108_/B VGND VPWR _1290_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_50_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_279 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1070_ _1070_/A _1070_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0923_ _0923_/X _2045_/Q _2044_/Q _2043_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1972_ _1972_/Q fanout174/X _1972_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1406_ _1406_/C _1406_/A _1407_/A _1406_/B _1405_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1268_ _1269_/B _1975_/Q _1267_/X _1266_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1337_ VGND VPWR _1436_/B _1337_/X _1429_/B _1729_/A VGND VPWR sky130_fd_sc_hd__and3b_2
X_1199_ VGND VPWR _1244_/A _1081_/Y _1198_/Y _1066_/A _1066_/C _1066_/D VGND VPWR
+ sky130_fd_sc_hd__a311o_2
XFILLER_43_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_117 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1122_ _1122_/C _1154_/A _1123_/D _1122_/B _1122_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_25_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1053_ _1160_/A _1053_/X _1090_/A _1053_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1886_ _2035_/D _1882_/Y _2035_/Q _1870_/C _1831_/B VGND VPWR _1885_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1955_ VGND VPWR _2063_/D _1955_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1671_ _1672_/B _1671_/C _2024_/Q _1671_/B _1671_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1740_ _2095_/A _1724_/A _1724_/B _1733_/A _1731_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_4
XFILLER_30_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xadc_core_digital_196 adc_core_digital_196/LO nmatrix_rowon_out_n[15] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
X_2085_ VGND VPWR _2085_/X _2085_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1105_ _1105_/B _1165_/A _1105_/A _1105_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1036_ _1036_/B _1036_/Y _1993_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1869_ VPWR VGND _1869_/X _1870_/C _2010_/Q _1870_/D _1869_/B VGND VPWR sky130_fd_sc_hd__and4b_2
X_1938_ VGND VPWR _2055_/D _1938_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1654_ _2021_/Q _1654_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1723_ _2084_/A _2081_/A _1744_/B _1712_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1585_ _1836_/A _2013_/Q _1584_/X _1585_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1019_ _1997_/Q _1157_/B _1995_/Q _1052_/C _1019_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_17_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_63 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1370_ _1469_/C _1370_/X _1731_/A _1457_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1637_ _1637_/Y _2018_/Q _1656_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1706_ VPWR VGND _1707_/A _1749_/B _1706_/D _1744_/B _2081_/A VGND VPWR sky130_fd_sc_hd__and4b_2
X_1568_ _1567_/X _1563_/X _2009_/Q _1665_/A _2009_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1499_ _1499_/Y _1977_/Q _2008_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_48_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1422_ _1422_/X _1413_/Y _1420_/Y _1419_/Y _1408_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1353_ _1353_/B _1353_/C _1353_/A _1353_/D _1354_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1284_ _1289_/B _1289_/A _1284_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
X_0999_ _2067_/Q input2/X _0999_/X _0998_/Y _2049_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_10_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0922_ _0921_/X _0919_/X _0916_/Y _0926_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1971_ _1971_/Q fanout175/X _1971_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1405_ _1405_/Y _1436_/B _1405_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1267_ VPWR VGND _1267_/A _1267_/X _1267_/B VGND VPWR sky130_fd_sc_hd__and2_2
Xinput1 VPWR VGND input1/X clk_dig_in VGND VPWR sky130_fd_sc_hd__buf_2
X_1336_ _1429_/B _1336_/A _1471_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1198_ _1198_/A _1198_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_19_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_97 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_272 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1121_ _1177_/B _1123_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1052_ _1052_/C _1053_/C _1995_/Q _1997_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_21_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1954_ VGND VPWR _1956_/D _1975_/D _1621_/A _1955_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1885_ _1884_/X _1883_/X _1923_/B _2016_/D _1885_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
XPHY_105 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1319_ _1355_/B _1320_/A _1471_/A _1412_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_8_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_95 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1670_ _1670_/B _2024_/D _1784_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_2084_ VGND VPWR _2084_/X _2084_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xadc_core_digital_197 adc_core_digital_197/LO pmatrix_c0_out_n VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__conb_1
X_1035_ VPWR VGND _1036_/B _1144_/A _1126_/A VGND VPWR sky130_fd_sc_hd__xor2_2
X_1104_ _1104_/A _1148_/A _1104_/C _1220_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
X_1937_ VGND VPWR _1977_/D _1967_/D _2055_/Q _1938_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1868_ _1513_/S _1867_/X _1866_/X _1868_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1799_ VGND VPWR _1799_/S _1997_/Q _1996_/Q _1800_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1653_ VPWR VGND _2018_/Q _1671_/C _2019_/Q VGND VPWR sky130_fd_sc_hd__and2_2
X_1722_ _2083_/A _1724_/A _1724_/B _1733_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_1584_ VGND VPWR _1584_/S _1579_/Y _2060_/Q _1584_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_2067_ _2067_/Q fanout175/X _2067_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1018_ VGND VPWR _1052_/C _1994_/Q _1996_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_17_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1705_ VPWR VGND _1744_/B _1729_/C VGND VPWR sky130_fd_sc_hd__buf_4
X_1567_ _1567_/A _1612_/B _2056_/Q _1567_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1636_ _1656_/B _1636_/X _2018_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1498_ _1498_/X _2055_/Q _1565_/A _1497_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_38_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1421_ _1421_/X _1418_/Y _1408_/A _1419_/Y _1420_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1352_ VPWR VGND _1353_/D _1352_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1283_ _1283_/C _1290_/A _1283_/X _1290_/B _1283_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0998_ _2067_/Q _0998_/Y _2066_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1619_ VPWR VGND _1619_/X _1619_/B _1606_/A VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_10_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1970_ _1970_/Q fanout178/X _1970_/D _2004_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_0921_ _0920_/Y _2046_/Q _0955_/B _0921_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_5_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1404_ _1404_/B _1406_/A _1435_/A _1404_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1335_ _1335_/X _1334_/X _1471_/A _1328_/Y _1305_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1197_ _1197_/B _1972_/D _1963_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xinput2 VPWR VGND input2/X comparator_in VGND VPWR sky130_fd_sc_hd__buf_4
X_1266_ _1245_/B _1266_/X _1265_/Y _1230_/X _1264_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o211a_4
XFILLER_2_284 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1051_ _1157_/B _1090_/A _1233_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1120_ _1119_/X _1262_/C _1157_/B _1187_/B _1154_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_4
X_1884_ _1915_/B _1884_/X _1928_/B _2014_/D _2012_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1953_ VGND VPWR _2062_/D _1953_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1318_ _1412_/B _1318_/A _1318_/B _1318_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_4
X_1249_ _1974_/D _1248_/Y _1259_/B _1717_/C _1963_/S _1717_/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a311oi_4
XPHY_106 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xadc_core_digital_198 adc_core_digital_198/LO pmatrix_rowon_out_n[15] VPWR VGND VGND
+ VPWR sky130_fd_sc_hd__conb_1
X_2083_ VGND VPWR _2083_/X _2083_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1034_ _2104_/A _1033_/Y _1216_/S _1966_/Q _1966_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1103_ _1103_/A _1104_/C _1103_/B _1103_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_2
X_1867_ _1928_/B _1867_/X _1867_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1936_ VGND VPWR _2054_/D _1936_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1798_ VGND VPWR _1995_/D _1798_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1721_ _2081_/A _1409_/B _2082_/A _1717_/B _1744_/B _1717_/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a41o_2
XFILLER_7_162 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1652_ _1671_/B _1634_/X _1606_/A _1632_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1583_ _2060_/Q _1893_/B _1583_/X _1582_/Y _1581_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_2066_ _2066_/Q fanout173/X _2066_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1017_ VGND VPWR _2005_/Q _1016_/X _1238_/C _1015_/Y _1014_/Y VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_34_283 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1919_ _1829_/B _1918_/X _1917_/Y _2021_/D _1919_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
XFILLER_17_217 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1704_ _1975_/Q _1729_/C _1269_/B _1267_/X _1266_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_2
X_1566_ VGND VPWR _1566_/S _1564_/Y _2009_/Q _1567_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1635_ _1634_/X _1632_/X _1606_/A _1656_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1497_ _1870_/A _1497_/Y _1496_/X _1621_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_2049_ _2049_/Q fanout175/X _2049_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_275 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1351_ VPWR VGND _1376_/A _1352_/A _1381_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1420_ _1706_/D _1420_/Y _1471_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_55_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1282_ _1289_/A _1289_/B _1283_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
X_1618_ VPWR VGND _1619_/B _1897_/C _1615_/Y VGND VPWR sky130_fd_sc_hd__and2b_2
X_0997_ VGND VPWR _0997_/S _0996_/X input2/X _0997_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1549_ _1612_/B _1552_/S _2014_/Q _1549_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_10_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0920_ _2065_/Q _0920_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_5_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1403_ _1403_/X _1405_/B _1332_/X _1406_/B _1406_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1265_ _1212_/B _1252_/X _1265_/Y _1222_/X _1212_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_2
X_1334_ _1334_/X _1460_/B _1706_/D _1469_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
Xinput3 VGND VPWR input3/X config_1_in[0] VGND VPWR sky130_fd_sc_hd__buf_1
X_1196_ VGND VPWR _1259_/B _1390_/A _1180_/B _1197_/B VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_296 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1050_ _1050_/A _1245_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_12
X_1883_ _2018_/D _1858_/A _1889_/B _1883_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1952_ VGND VPWR _1956_/D _1974_/D _2062_/Q _1953_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1248_ _1259_/B _1248_/Y _1974_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1317_ _1355_/B _1317_/A _1317_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_24_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1179_ VGND VPWR _1262_/B _1177_/X _1232_/B _1181_/B VGND VPWR sky130_fd_sc_hd__mux2_2
XPHY_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2082_ VGND VPWR _2082_/X _2082_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1102_ VGND VPWR _1993_/Q _1046_/A _1036_/B _1103_/C VGND VPWR sky130_fd_sc_hd__mux2_1
X_1033_ _1033_/Y _1216_/S _1033_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1866_ _1915_/A _2010_/Q _1866_/X _1870_/C _1928_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1935_ VGND VPWR _1977_/D _1966_/D _2054_/Q _1936_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1797_ VGND VPWR _1799_/S _1996_/Q _1995_/Q _1798_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_55 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1651_ _1651_/B _2020_/D _1784_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1720_ _2080_/A _1747_/B _1471_/B _1749_/D _1733_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_4
X_1582_ _2013_/Q _1582_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_19_281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_2065_ _2065_/Q fanout174/X _2065_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1016_ _1232_/B _2004_/Q _1232_/C _1016_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1849_ _1849_/X _1989_/Q _1849_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1918_ _1918_/X _1929_/S _2019_/Q _1917_/B _1882_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_48_321 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1634_ _1624_/X _1977_/Q _1633_/Y _1634_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1703_ _1749_/B _1717_/B _1717_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1565_ _1566_/S _1565_/A _1565_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1496_ _1500_/A _1496_/X _2008_/Q _1500_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_2048_ _2048_/Q fanout175/X _2048_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_13_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_98 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1350_ _1350_/B _1381_/B _1399_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1281_ _1281_/Y _1283_/C _1281_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_0_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0996_ _0996_/X _0995_/Y _2051_/Q _2065_/Q _2066_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1617_ _1897_/C _2063_/Q _2016_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1479_ _1984_/Q _1978_/Q _1480_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
X_1548_ _1543_/Y _1545_/X _1552_/S _1538_/C _1547_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_10_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_272 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1402_ _1402_/X _1397_/Y _1324_/X _1406_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
Xinput4 VGND VPWR input4/X config_1_in[1] VGND VPWR sky130_fd_sc_hd__buf_1
X_1264_ _1264_/Y _1264_/A _1264_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1333_ _1333_/X _1329_/Y _1332_/X _1328_/Y _1405_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_51_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1195_ _1318_/A _1318_/B _1318_/C _1390_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
X_0979_ _1233_/C _0980_/A _1122_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_10_58 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_99 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1882_ _1906_/A _1882_/Y _1882_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1951_ _2061_/D _1950_/X _1977_/D _2104_/A _1217_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1247_ _1246_/Y _1244_/Y _1245_/Y _1264_/A _1717_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_4
X_1178_ _1180_/B _1077_/D _1177_/X _1151_/X _0980_/A _1201_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_4
X_1316_ _1316_/A _1471_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
XPHY_108 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput160 VPWR VGND sample_switch_out _2105_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_127 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_2081_ VPWR VGND _2081_/X _2081_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1032_ _1032_/A _1033_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1101_ _1220_/A _1093_/X _1166_/A _1029_/X _1138_/A _1108_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
X_1934_ VGND VPWR _2053_/D _1934_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1865_ _1865_/X _1864_/Y _1893_/B _1864_/A _1870_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1796_ VGND VPWR _1994_/D _1796_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1650_ VGND VPWR _1651_/B _2020_/Q _1668_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1581_ VGND VPWR _1584_/S _2060_/Q _1579_/Y _1581_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_271 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1015_ _1015_/Y _1232_/C _2003_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_2064_ _2064_/Q fanout175/X _2064_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1917_ _1917_/Y _1929_/S _1917_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_1_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1779_ VPWR VGND _1780_/B _1779_/B _1986_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1848_ _1853_/A _1847_/X _1878_/B _1904_/A _1515_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1564_ _1564_/Y _1870_/A _2009_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1702_ VPWR VGND _2026_/D _1906_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1633_ _1633_/B _1633_/Y _1897_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1495_ _1621_/D _1906_/A _1697_/A _1478_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o21ai_4
X_2047_ _2047_/Q fanout174/X _2047_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_8_7 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1280_ _1289_/B _1281_/B _1289_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_51_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0995_ _2065_/Q _0994_/Y _2066_/Q _0995_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1616_ _2063_/Q _1626_/A _2016_/Q _1632_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1547_ _1547_/B _1547_/Y _1547_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1478_ _1981_/Q _1983_/Q _1979_/Q _1985_/Q _1478_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_54_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1401_ _1401_/X _1406_/C _1343_/A _1400_/X _1397_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1332_ VPWR VGND _1332_/X _1332_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xinput5 VGND VPWR input5/X config_1_in[2] VGND VPWR sky130_fd_sc_hd__buf_1
X_1263_ _1269_/A _1263_/B _1976_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
X_1194_ _1185_/X _1192_/Y _1318_/C _1190_/C _1193_/X _1191_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_0978_ _1151_/C _1233_/C _1157_/B _0978_/D _0990_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_15_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_180 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1950_ VPWR VGND _2061_/Q _1950_/X _1950_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1881_ _2034_/D _1877_/Y _1878_/X _1880_/X _1879_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1315_ _1315_/B _1316_/A _1315_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_24_114 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1246_ _1242_/A _1246_/Y _1245_/B _1973_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1177_ _2000_/Q _1999_/Q _1177_/X _1177_/B _2001_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
XFILLER_12_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput150 VPWR VGND result_out[2] _2029_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput161 VPWR VGND sample_switch_out_n _2106_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_294 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2080_ VGND VPWR _2080_/X _2080_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1100_ _1138_/A _1967_/Q _1099_/X _1041_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_38_206 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1031_ _1032_/A _1031_/B _1221_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1933_ VGND VPWR _1977_/D _1965_/D _2053_/Q _1934_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1864_ _1870_/B _1864_/Y _1864_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1795_ VGND VPWR _1799_/S _1995_/Q _1994_/Q _1796_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1229_ VGND VPWR _1201_/A _1229_/C _1227_/X _1229_/X _1229_/D VGND VPWR sky130_fd_sc_hd__and4bb_2
XFILLER_20_183 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_198 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_161 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1580_ _1537_/X _1539_/B _2012_/Q _1584_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_2063_ _2063_/Q fanout177/X _2063_/D _2063_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1014_ _2004_/Q _1014_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1847_ _1847_/B _1847_/X _2010_/Q _1878_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1916_ _1915_/X _1916_/Y _1861_/Y _1877_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1778_ _1779_/B _1985_/Q _1778_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_48_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1701_ _1819_/A _1906_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_31_289 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1563_ _1563_/X _2056_/Q _1507_/X _1562_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1632_ VGND VPWR _1632_/B _1632_/X _1633_/B _1977_/Q VGND VPWR sky130_fd_sc_hd__and3b_2
X_1494_ _1565_/A _2008_/Q _1500_/A _1500_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2046_ _2046_/Q fanout173/X _2046_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_1_138 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0994_ _2050_/Q _0994_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_5_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1477_ _1557_/B _2053_/Q _2006_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1615_ VGND VPWR _1615_/Y _2064_/Q _2017_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1546_ VGND VPWR _1547_/B _2012_/Q _2059_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_42_318 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_2029_ _2029_/Q fanout165/X _2029_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_18_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1331_ _1436_/B _1332_/A _1435_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1400_ _1469_/C _1400_/X _1469_/A _1460_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1262_ _1262_/B _1262_/C _1262_/A _1262_/D _1263_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
X_1193_ _1193_/B _1193_/X _1193_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_36_101 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput6 VPWR VGND input6/X config_1_in[3] VGND VPWR sky130_fd_sc_hd__buf_2
X_0977_ _2105_/A _1992_/Q _0978_/D _1993_/Q _1991_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
XFILLER_19_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1529_ _1529_/A _1529_/B _1529_/C _1538_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_35_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_23 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_266 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_134 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1880_ _1906_/C _1880_/X _1861_/Y _2034_/Q _2056_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_18_189 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_90 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_192 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1314_ _1314_/Y _1469_/A _1469_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_4
X_1245_ _1245_/Y _1973_/Q _1245_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_49_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1176_ VGND VPWR _1262_/C _1227_/B _1193_/B _1151_/X _1150_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_21_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput151 VPWR VGND result_out[3] _2030_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput140 VPWR VGND pmatrix_rowon_out_n[8] _2097_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1030_ _1220_/A _1029_/X _1031_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2b_2
X_1932_ _2042_/D _1931_/X _1930_/X _1858_/A _1928_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1863_ _1856_/Y _1862_/X _1860_/X _2032_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1794_ VGND VPWR _1993_/D _1794_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1228_ VGND VPWR _1232_/B _1160_/A _1057_/Y _1229_/C VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1159_ VGND VPWR _1155_/X _1245_/B _1187_/B _1166_/B _1158_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_2062_ _2062_/Q fanout177/X _2062_/D _2063_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1013_ VPWR VGND _1262_/B _1151_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1777_ _1777_/B _1985_/D _2026_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1846_ _1920_/B _1878_/B _1929_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1915_ _1915_/C _1915_/A _1915_/X _1915_/B _1915_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_25_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1700_ _1819_/A _1882_/A _1751_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1631_ VPWR VGND _2017_/D _1631_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_31_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1562_ _1864_/A _1562_/Y _1508_/X _1612_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1493_ _1500_/B _2054_/Q _2006_/Q _2007_/Q _2053_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_2045_ _2045_/Q fanout173/X _2045_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_224 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1829_ VPWR VGND _1917_/B _1833_/B _1829_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_13_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_239 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0993_ _0993_/A _1007_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1614_ VPWR VGND _2016_/D _1614_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1476_ VPWR VGND _1882_/A _1836_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1545_ _1545_/X _2013_/Q _2012_/Q _2060_/Q _2059_/Q VGND VPWR _1544_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_2028_ _2028_/Q fanout165/X _2028_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_49_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1261_ _2005_/Q _1262_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1330_ _1330_/X _1324_/X _1405_/B _1328_/Y _1329_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
Xinput7 VPWR VGND input7/X config_1_in[4] VGND VPWR sky130_fd_sc_hd__buf_2
X_1192_ _1192_/Y _1193_/A _1193_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0976_ VPWR VGND _1233_/C _1122_/D VGND VPWR sky130_fd_sc_hd__buf_6
X_1528_ _1529_/C _1500_/A _2054_/Q _1526_/X _1527_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1459_ _1459_/X _1452_/Y _1451_/B _1427_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_51_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1244_ _1244_/Y _1244_/A _1244_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_49_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1313_ VPWR VGND _1469_/C _1436_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1175_ _1971_/Q _1227_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_0959_ _1965_/Q _1145_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
Xoutput141 VPWR VGND pmatrix_rowon_out_n[9] _2098_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput152 VPWR VGND result_out[4] _2031_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput130 VPWR VGND pmatrix_rowon_out_n[12] _2101_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_46_285 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1931_ _2042_/Q _1819_/A _1931_/X _2017_/D _1882_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1862_ _1906_/C _1862_/X _1861_/Y _2032_/Q _2007_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1793_ VGND VPWR _1793_/S _1994_/Q _1993_/Q _1794_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1227_ _1232_/C _1227_/B _1227_/X _1227_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1158_ _1158_/A _1158_/B _1158_/X _1158_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1089_ VPWR VGND _1090_/B _1157_/C _1156_/A _1089_/C _1156_/B VGND VPWR sky130_fd_sc_hd__and4b_2
XFILLER_28_230 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_277 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_241 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_2061_ _2061_/Q fanout175/X _2061_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1012_ _1966_/Q _1065_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1914_ VGND VPWR _1915_/D _2019_/Q _1914_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1845_ _2030_/Q _1831_/B _2030_/D _1844_/X _1842_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1776_ VGND VPWR _1777_/B _1985_/Q _1778_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_25_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_288 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1630_ VGND VPWR _1631_/A _1629_/X _1622_/Y _1665_/A _1869_/B _1620_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_2
X_1561_ _1558_/Y _2007_/Q _2007_/D _1893_/B _1560_/X _1665_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1492_ _1500_/A _2007_/Q _2053_/Q _2006_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2044_ _2044_/Q fanout173/X _2044_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1759_ _1760_/S _1978_/Q _1979_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1828_ VGND VPWR _1929_/S _2010_/D _2008_/D _1828_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0992_ _1221_/B _0993_/A _0992_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1613_ _1621_/A _1893_/A _1614_/A _1608_/X _1612_/X _1665_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1544_ _1519_/B _1524_/A _2059_/Q _2012_/Q _1544_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1475_ _1596_/A _1836_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
X_2027_ _2027_/Q fanout165/X _2027_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_42_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xinput8 VPWR VGND input8/X config_1_in[5] VGND VPWR sky130_fd_sc_hd__buf_2
X_1191_ _1203_/B _1191_/Y _1203_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1260_ _1258_/Y _2104_/A _1259_/X _1975_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_36_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0975_ _1997_/Q _1994_/Q _1122_/D _1995_/Q _1996_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_10_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1527_ _2056_/Q _2009_/Q _1527_/X _2008_/Q _2055_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1389_ _1749_/A _1391_/A _1435_/B _1404_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_27_136 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1458_ _1458_/X _1451_/B _1343_/A _1454_/X _1457_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_50_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1312_ VPWR VGND _1436_/B _1349_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1243_ _1242_/X _1219_/Y _1231_/X _1973_/Q _1717_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_4
X_1174_ _1029_/X _1138_/A _1093_/X _1220_/A _1190_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_0958_ _0958_/B _2047_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xoutput142 VPWR VGND result_out[0] _2027_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput120 VPWR VGND pmatrix_row_out_n[3] _2091_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput131 VPWR VGND pmatrix_rowon_out_n[13] _2102_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput153 VPWR VGND result_out[5] _2032_/Q VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1930_ _1889_/B _1930_/X _1929_/X _2025_/D _1920_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_46_297 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1861_ _1861_/Y _1904_/A _1861_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1792_ VGND VPWR _1992_/D _1792_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1157_ _1157_/C _1233_/A _1158_/C _1157_/B _1089_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1226_ _1226_/B _1226_/Y _1226_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1088_ VPWR VGND _1089_/C _1126_/A _1997_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_7_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2060_ _2060_/Q fanout168/X _2060_/D _2060_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1011_ _2104_/A _1007_/Y _1216_/S _1965_/Q _1965_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1913_ _1913_/B _1914_/B _1913_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1844_ _1889_/B _1844_/X _2013_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1775_ _1984_/Q _1778_/B _1983_/Q _1775_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_25_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1209_ _1344_/B _1208_/Y _1244_/A _1244_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_40_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1560_ _1560_/X _2054_/Q _1500_/A _1559_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1491_ VPWR VGND _1864_/A _1870_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_2043_ _2043_/Q _2043_/D VPWR fanout173/X _2066_/CLK VGND VGND VPWR sky130_fd_sc_hd__dfstp_4
X_1827_ _2028_/D _1826_/X _1825_/X _2026_/D _1822_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1758_ _1882_/A _1758_/Y _1980_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1689_ _1920_/B _1690_/A _1987_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_45_307 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_292 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_81 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_178 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_270 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0991_ _1221_/B _1145_/A _1105_/B _0990_/D _0990_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_4
X_1612_ _1612_/A _1612_/B _1621_/A _1612_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1474_ _1977_/Q _1596_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1543_ _1547_/A _1543_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_2026_ _2026_/Q fanout169/X _2026_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput9 VGND VPWR input9/X rst_n VGND VPWR sky130_fd_sc_hd__buf_1
X_1190_ _1190_/A _1190_/B _1318_/B _1190_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_0974_ _0968_/X _0965_/X _1105_/B _1223_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
X_1526_ _2053_/Q _1526_/X _2007_/Q _2006_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1457_ _1469_/C _1457_/X _1464_/A _1457_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1388_ VGND VPWR _1388_/X _1388_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_2009_ _2009_/Q fanout165/X _2009_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_14_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1311_ VPWR VGND _1311_/A _1349_/C _1311_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_1_291 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1242_ _1242_/A _1242_/B _1241_/X _1242_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1173_ _1220_/B _1173_/B _1190_/A _1173_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
Xoutput121 VPWR VGND pmatrix_row_out_n[4] _2092_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput110 VPWR VGND pmatrix_col_out_n[8] _1347_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_0957_ VPWR VGND _0958_/B _0957_/B _2047_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
Xoutput132 VPWR VGND pmatrix_rowon_out_n[14] _2103_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput143 VPWR VGND result_out[10] _2037_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput154 VPWR VGND result_out[6] _2033_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1509_ _1508_/X _1507_/X _2056_/Q _1513_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_55_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1860_ _1860_/X _1906_/D _2013_/D _1857_/Y _1859_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1791_ VGND VPWR _1793_/S _1993_/Q _1992_/Q _1792_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1087_ VGND VPWR _1968_/D _1087_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_257 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1156_ _1158_/B _1156_/A _1156_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1225_ VGND VPWR _1267_/A _1224_/Y _1198_/Y _1066_/C _1220_/Y _1221_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_2
X_1989_ _1989_/Q fanout166/X _1989_/D _2039_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_4_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1010_ VGND VPWR _2106_/A _1956_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_1843_ _1889_/B _1989_/Q _1849_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_1912_ _1909_/X _1911_/X _1910_/X _2039_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1774_ _1774_/B _1984_/D _2026_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1208_ _1208_/Y _1289_/B _1290_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1139_ _1138_/C _1315_/B _1138_/D _1138_/Y _1211_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22ai_4
X_1490_ _1882_/A _1489_/X _1485_/X _2006_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_2042_ _2042_/Q fanout170/X _2042_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_249 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1826_ VPWR VGND _2028_/Q _1826_/X _1831_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1757_ _1756_/X _1979_/D _1755_/X _1754_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1688_ _1988_/Q _1989_/Q _1920_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2b_4
XFILLER_45_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_71 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_282 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1611_ VGND VPWR _1897_/A _1893_/A _1610_/Y _1612_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_0990_ _0992_/A _0990_/C _1145_/A _1105_/B _0990_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1542_ _2060_/Q _1547_/A _2013_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1473_ _1473_/X _1451_/A _1412_/Y _1409_/B _1314_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_2025_ _2025_/Q fanout169/X _2025_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_54_127 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1809_ VGND VPWR _1817_/S _1232_/C _1126_/A _1810_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0973_ _1223_/A _1233_/A _1157_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1525_ _1529_/B _2009_/Q _2056_/Q _2055_/Q _2008_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1387_ _1391_/C _1387_/A _1388_/A _1391_/B _1386_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1456_ _1456_/X _1368_/Y _1408_/B _1446_/X _1454_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_23_322 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2008_ _2008_/Q fanout167/X _2008_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_50_163 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_237 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_281 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1310_ _1309_/Y _1307_/Y _1305_/X _1409_/B _1310_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1241_ _1290_/B _1212_/A _1238_/X _1290_/A _1241_/X _1212_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_1172_ _1180_/B _1972_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_49_252 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0956_ _0956_/B _2046_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xoutput100 VPWR VGND pmatrix_col_out_n[28] _1403_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput111 VPWR VGND pmatrix_col_out_n[9] _1354_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput155 VPWR VGND result_out[7] _2034_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput122 VPWR VGND pmatrix_row_out_n[5] _2093_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput144 VPWR VGND result_out[11] _2038_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput133 VPWR VGND pmatrix_rowon_out_n[1] _2090_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1508_ _1565_/A _1508_/X _2009_/Q _1565_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1439_ _1439_/X _1367_/X _1413_/Y _1368_/Y _1430_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_23_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_174 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1790_ VGND VPWR _1991_/D _1790_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1224_ _1223_/X _1104_/A _1224_/Y _1104_/C _1222_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a31oi_2
X_1086_ VPWR VGND _1956_/B _1087_/A _1086_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_52_269 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1155_ _1123_/D _1119_/X _1154_/X _1238_/C _1020_/X _1155_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_1988_ _1988_/Q fanout165/X _1988_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0939_ input2/X _0942_/B _2048_/Q _2049_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_43_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_95 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout190 VPWR VGND _2005_/CLK _2063_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1773_ VPWR VGND _1774_/B _1773_/B _1984_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
X_1842_ _1920_/B _1835_/X _1842_/X _1837_/X _1841_/X _1923_/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1911_ _1906_/C _1911_/X _1861_/Y _2039_/Q _2061_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1207_ _1290_/C _1212_/A _1206_/X _1203_/B _1203_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_4
XFILLER_25_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1138_ _1166_/A _1138_/A _1138_/Y _1138_/D _1138_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4_2
X_1069_ VPWR VGND _1070_/A _1069_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_324 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2041_ _2041_/Q fanout170/X _2041_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_54_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1756_ _1979_/Q _1756_/B _1978_/Q _1756_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1825_ _2011_/D _1920_/B _1825_/X _2009_/D _1906_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1687_ _1686_/X _1904_/C _1682_/X _1989_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_36_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1610_ _1610_/Y _1870_/A _2016_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1541_ _2012_/D _1850_/B _1850_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1472_ _1471_/Y _1405_/Y _1464_/X _1409_/B _1472_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_2024_ _2024_/Q fanout171/X _2024_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1808_ VGND VPWR _2000_/D _1808_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1739_ _1733_/A _1724_/B _1724_/A _2094_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_14_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_93 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0972_ VPWR VGND _1157_/B _1122_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1524_ _1529_/A _1867_/A _1524_/A _1524_/B _1524_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1386_ _1386_/Y _1436_/B _1386_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1455_ _1455_/X _1454_/X _1413_/Y _1368_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2007_ _2007_/Q fanout167/X _2007_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_14_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1171_ _2104_/A _1170_/Y _1216_/S _1971_/Q _1971_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1240_ _1173_/B _1138_/A _1166_/A _1220_/B _1290_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_4
X_0955_ VGND VPWR _0956_/B _2046_/Q _0955_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
Xoutput145 VPWR VGND result_out[12] _2039_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput134 VPWR VGND pmatrix_rowon_out_n[2] _2091_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput101 VPWR VGND pmatrix_col_out_n[29] _1407_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1507_ _1507_/X _2009_/Q _1565_/A _1565_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
Xoutput123 VPWR VGND pmatrix_row_out_n[6] _2094_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput156 VPWR VGND result_out[8] _2035_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput112 VPWR VGND pmatrix_row_out_n[10] _2098_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1369_ _1408_/B _1368_/Y _1359_/C _1366_/X _1367_/X _1369_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a221oi_2
X_1438_ _1438_/X _1433_/X _1314_/Y _1368_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_46_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1223_ _1223_/A _1262_/B _1053_/C _1223_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1154_ _1233_/C _1154_/X _1154_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1085_ VGND VPWR _1259_/B _1435_/A _1968_/Q _1086_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_1987_ _1987_/Q fanout165/X _1987_/D _2034_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0938_ _0938_/B _2049_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_51_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout180 VPWR VGND _2039_/CLK fanout186/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_256 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout191 VPWR VGND _2063_/CLK _2004_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
X_1910_ _1910_/X _1849_/X _2016_/D _2022_/D _1870_/D VGND VPWR _1915_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1772_ _1773_/B _1983_/Q _1775_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1841_ _1858_/A _1839_/X _1928_/B _2007_/D _1841_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1206_ _1206_/X _1155_/X _1138_/D _1201_/A _1201_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1137_ VGND VPWR _1136_/Y _1211_/B _1165_/C _1131_/Y _1315_/A _1135_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_4
X_1068_ VPWR VGND _1069_/A _1068_/B _1066_/X VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_48_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_130 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_2040_ _2040_/Q fanout170/X _2040_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_15_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1755_ _1755_/X _1978_/Q _1861_/B _1904_/A _1840_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1686_ _1829_/B _1984_/Q _1686_/X _1686_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1824_ _1917_/B _1906_/D _1929_/S _1829_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_38_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_177 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_115 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1540_ _1539_/Y _1537_/X _1836_/A _1850_/C _2012_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_4
XFILLER_10_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1471_ _1471_/Y _1471_/A _1471_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_2023_ _2023_/Q fanout169/X _2023_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1807_ VGND VPWR _1817_/S _1126_/A _1144_/A _1808_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1669_ _1670_/B _1669_/B _2024_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xor2_4
X_1738_ _2081_/A _1712_/C _1744_/B _2093_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_14_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0971_ _2003_/Q _2005_/Q _1122_/C _2004_/Q _2002_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XFILLER_4_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1523_ _2057_/Q _1524_/D _2056_/Q _2010_/Q _2009_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1454_ _1454_/X _1451_/B _1464_/A _1399_/A _1729_/A VGND VPWR _1394_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1385_ _1385_/X _1386_/B _1332_/X _1391_/B _1391_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_2006_ _2006_/Q fanout167/X _2006_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1170_ _1170_/Y _1216_/S _1350_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0954_ _0954_/B _2045_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xoutput102 VPWR VGND pmatrix_col_out_n[2] _1322_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput135 VPWR VGND pmatrix_rowon_out_n[3] _2092_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1506_ _1565_/B _2055_/Q _1500_/B _2008_/Q _1500_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
Xoutput157 VPWR VGND result_out[9] _2036_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput146 VPWR VGND result_out[13] _2040_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput113 VPWR VGND pmatrix_row_out_n[11] _2099_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput124 VPWR VGND pmatrix_row_out_n[7] _2095_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1437_ _1437_/X _1368_/Y _1343_/A _1433_/X _1436_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1299_ VPWR VGND _1706_/D _1729_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1368_ _1368_/Y _1471_/A _1412_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_11_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1153_ VGND VPWR _1162_/B _1971_/Q _1188_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1222_ _1262_/B _1222_/X _1262_/C _1238_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or3_4
X_1084_ VPWR VGND _1435_/A _1336_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1986_ _1986_/Q fanout169/X _1986_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0937_ VPWR VGND _0938_/B _0937_/B _2049_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_28_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_146 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout170 VPWR VGND fanout170/X fanout171/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout181 VPWR VGND _2059_/CLK fanout186/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout192 VPWR VGND _2004_/CLK input1/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_61 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1840_ _1864_/A _1906_/A _1840_/C _1858_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
X_1771_ _1771_/B _1983_/D _2026_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1067_ _1066_/A _1081_/A _1068_/B _1066_/D _1066_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1136_ _1173_/B _1138_/C _1173_/C _1166_/A _1138_/A _1136_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a2111oi_4
X_1205_ _1289_/B _1245_/B _1973_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1969_ _1969_/Q fanout173/X _1969_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1823_ _2027_/Q _1831_/B _2027_/D _2010_/D _1822_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_15_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1754_ _1979_/Q _1754_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1685_ VGND VPWR _1686_/C _1978_/Q _1849_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_2099_ VGND VPWR _2099_/X _2099_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1119_ _1119_/X _1117_/Y _1156_/A _1118_/X _1123_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_28_63 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_245 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1470_ _1731_/A _1405_/B _1408_/Y _1470_/Y _1469_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_2
X_2022_ _2022_/Q fanout169/X _2022_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1806_ VGND VPWR _1999_/D _1806_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1668_ _1669_/B _1668_/A _1671_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1599_ VPWR VGND _1877_/A _1599_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1737_ _1744_/B _2092_/A _2081_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_26_322 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0970_ VPWR VGND _1233_/A _1122_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1522_ _1867_/A _2010_/Q _2057_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1453_ _1453_/X _1451_/X _1314_/Y _1452_/Y _1368_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1384_ _1384_/X _1391_/B _1324_/X _1391_/C _1386_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_2005_ _2005_/Q fanout176/X _2005_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_64 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_97 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput114 VPWR VGND pmatrix_row_out_n[12] _2100_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput125 VPWR VGND pmatrix_row_out_n[8] _1724_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_0953_ VPWR VGND _0954_/B _0953_/B _2045_/Q VGND VPWR sky130_fd_sc_hd__xor2_2
Xoutput103 VPWR VGND pmatrix_col_out_n[30] _1410_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput158 VPWR VGND sample_matrix_out _2105_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput136 VPWR VGND pmatrix_rowon_out_n[4] _2093_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1505_ _1621_/D _1505_/Y _1870_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xoutput147 VPWR VGND result_out[14] _2041_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1367_ VPWR VGND _1399_/A _1367_/X _1367_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1436_ _1436_/B _1436_/X _1749_/A _1464_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1298_ VPWR VGND _1729_/A _1376_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_11_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_166 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1221_ _1221_/B _1221_/X _1966_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1152_ _1151_/X _1150_/X _1188_/B _0980_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_4
X_1083_ _1336_/A _1083_/B _1083_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
X_1985_ _1985_/Q fanout169/X _1985_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0936_ _0937_/B _2048_/Q input2/X VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1419_ _1460_/B _1419_/Y _1706_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_51_250 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout182 VPWR VGND _2060_/CLK fanout186/X VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout171 VPWR VGND fanout171/X fanout172/X VGND VPWR sky130_fd_sc_hd__buf_6
X_1770_ VGND VPWR _1771_/B _1983_/Q _1775_/C VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_6_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1204_ _1173_/B _1212_/B _1212_/A _1244_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1066_ _1066_/X _1066_/C _1066_/A _1081_/A _1066_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1135_ _1138_/D _1138_/C _1173_/C _1173_/B _1135_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1899_ _2014_/D _1898_/X _1928_/B _1899_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1968_ _1968_/Q fanout174/X _1968_/D _2065_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0919_ _0919_/X _0918_/X _0917_/X _2046_/Q _2045_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_0_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_86 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1753_ VGND VPWR _1978_/D _1753_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1822_ _1906_/C _1822_/X _1920_/B _1822_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1684_ _1849_/B _1987_/Q _1988_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_2098_ VGND VPWR _2098_/X _2098_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1118_ _1177_/B _1144_/A _1126_/A _1118_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1049_ _1229_/D _1050_/A _1160_/A _1160_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_0_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2021_ _2021_/Q fanout169/X _2021_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_39_128 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1736_ VGND VPWR _2091_/A _1736_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1805_ VGND VPWR _1817_/S _1144_/A _1123_/A _1806_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1667_ _1671_/D _2022_/Q _2020_/Q _2021_/Q _2023_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1598_ VPWR VGND _1599_/A _1588_/X _1598_/D _1598_/C _1598_/B VGND VPWR sky130_fd_sc_hd__and4b_2
X_1521_ _1524_/B _2011_/Q _1836_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1383_ _1451_/B _1391_/C _1464_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1452_ _1412_/B _1731_/A _1435_/B _1452_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_2004_ _2004_/Q fanout178/X _2004_/D _2004_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_50_112 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1719_ _1747_/B _1724_/B _1733_/A _2079_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_18_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_252 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_0952_ _0953_/B _2044_/Q _2043_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_32_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput159 VPWR VGND sample_matrix_out_n _2104_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput115 VPWR VGND pmatrix_row_out_n[13] _2101_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput126 VPWR VGND pmatrix_row_out_n[9] _2097_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1504_ VPWR VGND _1870_/C _2057_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput104 VPWR VGND pmatrix_col_out_n[31] _1411_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput148 VPWR VGND result_out[15] _2042_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput137 VPWR VGND pmatrix_rowon_out_n[5] _2094_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1435_ _1435_/B _1464_/C _1435_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1366_ VPWR VGND _1366_/X _1464_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1297_ _1376_/A _1344_/B _1344_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_55_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1220_ _1220_/B _1220_/Y _1220_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1151_ _1232_/B _1227_/C _1151_/C _1232_/C _1151_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__or4b_4
X_1082_ _1083_/B _1081_/Y _1066_/D _1066_/A _1066_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1984_ _1984_/Q fanout169/X _1984_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0935_ VPWR VGND _1799_/S _1817_/S VGND VPWR sky130_fd_sc_hd__buf_6
X_1349_ _1376_/A _1353_/C _1435_/B _1349_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1418_ _1408_/B _1418_/Y _1731_/A _1469_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_51_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout183 VPWR VGND _2026_/CLK _2024_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout172 VPWR VGND fanout172/X input9/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_8_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1134_ _1158_/A _1223_/A _1090_/B _1138_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__or3b_4
X_1203_ _1202_/X _1203_/B _1226_/A _1203_/A _1212_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or4b_4
XFILLER_18_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1065_ _1066_/D _1065_/A _1065_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1898_ _1906_/A _1897_/X _1896_/X _1915_/B _1898_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_0918_ _2066_/Q _2067_/Q _2065_/Q _0918_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1967_ _1967_/Q fanout173/X _1967_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_33_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1752_ VGND VPWR _1978_/Q _1756_/B _1904_/A _1753_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1683_ _1989_/Q _1829_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1821_ _1870_/D _1822_/C _1861_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_2097_ VGND VPWR _2097_/X _2097_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1117_ VGND VPWR _1117_/Y _1177_/B _1126_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1048_ _1015_/Y _2005_/Q _1016_/X _1160_/C _1014_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a211oi_2
XFILLER_0_158 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2020_ _2020_/Q fanout171/X _2020_/D _2024_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1666_ _1663_/Y _1786_/S _1664_/X _2023_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1735_ _1749_/D _1736_/A _1747_/B _1735_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1804_ VGND VPWR _1998_/D _1804_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1597_ VGND VPWR _1597_/S _1596_/X _1595_/X _1598_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1520_ VPWR VGND _1836_/C _2058_/Q VGND VPWR sky130_fd_sc_hd__buf_4
X_1451_ VPWR VGND _1451_/A _1451_/X _1451_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1382_ VPWR VGND _1391_/B _1382_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_2003_ _2003_/Q fanout178/X _2003_/D _2004_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1649_ _1656_/C _1668_/A _1656_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1718_ _1724_/A _1735_/C _1724_/B _2078_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_187 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_0951_ _0951_/B _2044_/D _1799_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_32_124 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput116 VPWR VGND pmatrix_row_out_n[14] _2102_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput149 VPWR VGND result_out[1] _2028_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput127 VPWR VGND pmatrix_rowon_out_n[0] _2089_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1503_ _1502_/X _1498_/X _2008_/Q _1864_/A _2008_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
Xoutput105 VPWR VGND pmatrix_col_out_n[3] _1330_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput138 VPWR VGND pmatrix_rowon_out_n[6] _2095_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1296_ _1471_/B _1423_/B _1408_/A _1296_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1365_ _1365_/X _1364_/X _1412_/B _1363_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1434_ _1434_/X _1367_/B _1408_/B _1432_/X _1433_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_11_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1150_ _1157_/B _1150_/B _1150_/X _1150_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1081_ _1081_/A _1081_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1983_ _1983_/Q fanout169/X _1983_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0934_ VPWR VGND _1817_/S _0934_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1417_ _1409_/B _1416_/X _1405_/B _1309_/Y _1417_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_4
X_1348_ _1429_/B _1353_/B _1464_/A _1436_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor3_2
X_1279_ _1226_/A _1203_/B _1203_/A _1283_/C _1212_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_4
XFILLER_51_274 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xfanout184 VPWR VGND _2042_/CLK _2024_/CLK VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_216 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout162 _2096_/A _1724_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout173 VPWR VGND fanout173/X fanout174/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_6_186 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1202_ _1969_/Q _1202_/B _1155_/X _1202_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_1133_ _1969_/Q _1158_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1064_ _1148_/A _1148_/B _1065_/B _1114_/D _1148_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_18_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1966_ _1966_/Q fanout173/X _1966_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1897_ _1897_/C _1897_/A _1897_/X _1915_/A _1915_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_0917_ _2043_/Q _0917_/X _2044_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1820_ _1917_/B _1870_/D _1987_/Q _1829_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_15_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1751_ _1756_/B _1904_/A _1751_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1682_ _1681_/Y _1978_/Q _1480_/D _1917_/B _1987_/Q _1682_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
X_1047_ _1233_/C _1229_/D _1233_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1116_ _1220_/B _1211_/B _1065_/B _1114_/X _1115_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22ai_4
X_2096_ VGND VPWR _2096_/X _2096_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_266 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1949_ _1956_/D _1950_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_44_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_185 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1803_ VGND VPWR _1817_/S _1123_/A _1177_/B _1804_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1665_ _1786_/S _1665_/A _1893_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1596_ _2015_/Q _1596_/A _1596_/X _2062_/Q _1621_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1734_ VPWR VGND _2090_/A _1734_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_2079_ VGND VPWR _2079_/X _2079_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_89 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1450_ _1450_/Y _1324_/X _1449_/X _1391_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21boi_4
X_1381_ VPWR VGND _1404_/B _1382_/A _1381_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_2002_ _2002_/Q fanout178/X _2002_/D _2004_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_35_144 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1648_ _1656_/C _2018_/Q _2019_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1579_ _1612_/B _1579_/Y _2060_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1717_ _1735_/C _1729_/A _1717_/B _1717_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand3_4
XPHY_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_0950_ VGND VPWR _0951_/B _2044_/Q _2043_/Q VGND VPWR sky130_fd_sc_hd__xnor2_2
Xoutput117 VPWR VGND pmatrix_row_out_n[15] _2103_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput128 VPWR VGND pmatrix_rowon_out_n[10] _2099_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1502_ _1502_/A _1621_/D _2055_/Q _1502_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
Xoutput106 VPWR VGND pmatrix_col_out_n[4] _1333_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput139 VPWR VGND pmatrix_rowon_out_n[7] _2096_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_49_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1433_ _1433_/X _1367_/B _1464_/A _1399_/A _1749_/A VGND VPWR _1423_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1364_ _1364_/X _1386_/B _1381_/B _1729_/A _1436_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1295_ VPWR VGND _1471_/B _1731_/A VGND VPWR sky130_fd_sc_hd__buf_6
X_1080_ _1083_/A _1211_/A _1198_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1982_ _1982_/Q fanout169/X _1982_/D _2026_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0933_ VGND VPWR _2048_/D input2/X _0933_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1347_ _1347_/X _1353_/A _1343_/Y _1435_/B _1409_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1416_ _1435_/A _1706_/D _1416_/X _1446_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1278_ VPWR VGND _1408_/A _1278_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_3_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout185 VPWR VGND _2024_/CLK fanout186/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout163 VPWR VGND _2081_/A _1271_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout174 VPWR VGND fanout174/X fanout177/X VGND VPWR sky130_fd_sc_hd__buf_6
X_1201_ _1226_/A _1201_/A _1201_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1063_ _0990_/C _1114_/D _0989_/B _1145_/A _1062_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1132_ _1245_/B _1138_/C _1129_/X _1187_/B _1123_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o211a_4
X_0916_ _0916_/Y _2066_/Q _0997_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1965_ _1965_/Q fanout175/X _1965_/D _2067_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1896_ _1893_/A _1896_/X _1786_/S _1904_/A _1621_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
XFILLER_3_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_179 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1750_ VPWR VGND _2103_/A _1750_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1681_ _1680_/X _1679_/Y _1987_/Q _1681_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_2_190 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_2095_ VGND VPWR _2095_/X _2095_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1046_ VPWR VGND _1046_/A _1160_/A _1156_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1115_ _1115_/X _1065_/A _1104_/C _1104_/A _1148_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1879_ _1879_/X _1849_/X _2011_/D _2017_/D _1870_/D VGND VPWR _1915_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_21_234 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1948_ VGND VPWR _2060_/D _1948_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1733_ _1747_/B _1734_/A _1733_/A _1749_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1802_ VGND VPWR _1997_/D _1802_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1664_ _1671_/B _1664_/X _1664_/A _1664_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1595_ _1596_/A _2015_/Q _2062_/Q _1595_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
X_2078_ VGND VPWR _2078_/X _2078_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1029_ _1029_/X _1065_/A _1148_/A _1148_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_55_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1380_ _1380_/X _1379_/X _1412_/B _1378_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2001_ _2001_/Q fanout178/X _2001_/D _2004_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_50_137 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1716_ _1724_/B _2077_/A _1724_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1578_ _1869_/B _1570_/Y _2011_/D _1836_/B _1904_/A _1857_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221ai_2
X_1647_ _2019_/D _1646_/X _2019_/Q _1643_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XPHY_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_167 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_299 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput107 VPWR VGND pmatrix_col_out_n[5] _1335_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_40_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1501_ VGND VPWR _1501_/S _1499_/Y _2008_/Q _1502_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput118 VPWR VGND pmatrix_row_out_n[1] _2089_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput129 VPWR VGND pmatrix_rowon_out_n[11] _2100_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1432_ _1446_/B _1432_/X _1464_/A _1457_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1363_ _1367_/B _1446_/B _1363_/X _1469_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
X_1294_ VPWR VGND _1731_/A _1749_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_11_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_284 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_89 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1981_ _1981_/Q fanout170/X _1981_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0932_ _0933_/B _2048_/Q _0949_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_45_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1346_ _1367_/B _1353_/A _1464_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1415_ _1415_/X _1321_/Y _1408_/A _1423_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1277_ _1350_/B _1278_/A _1399_/A _1464_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
Xfanout186 VPWR VGND fanout186/X input1/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_262 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xfanout164 VPWR VGND _2104_/A _2106_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout175 VPWR VGND fanout175/X fanout177/X VGND VPWR sky130_fd_sc_hd__buf_6
X_1200_ _1201_/B _1201_/A _1193_/B _1212_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ba_4
X_1062_ _1145_/A _1233_/A _1062_/X _1233_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1131_ _1289_/A _1131_/Y _1173_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_33_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1895_ _1923_/B _1895_/X _1894_/X _2018_/D _1915_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1964_ VGND VPWR _2067_/D _1964_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0915_ _2067_/Q _0997_/S VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_33_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_265 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1329_ _1731_/A _1329_/Y _1451_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_33_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1680_ VGND VPWR _1987_/Q _1982_/Q _1984_/Q _1680_/X _1988_/Q VGND VPWR sky130_fd_sc_hd__and4bb_2
XFILLER_24_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1114_ _1114_/X _1148_/D _1148_/A _1148_/B _1114_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1045_ _1144_/A _1046_/A _1126_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_2094_ VGND VPWR _2094_/X _2094_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1878_ VPWR VGND _2013_/D _1878_/X _1878_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1947_ VGND VPWR _1956_/D _1972_/D _2060_/Q _1948_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1663_ _1664_/A _1664_/C _1671_/B _1663_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1732_ VPWR VGND _2089_/A _1732_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1801_ VGND VPWR _1817_/S _1177_/B _1997_/Q _1802_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1594_ VGND VPWR _1597_/S _1605_/A _1590_/X _1598_/C VGND VPWR sky130_fd_sc_hd__mux2_1
X_2077_ VGND VPWR _2077_/X _2077_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_305 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1028_ _1065_/A _1148_/A _1148_/B _1220_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_17_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2000_ _2000_/Q fanout176/X _2000_/D _2005_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1646_ _1913_/A _1645_/Y _1913_/B _1646_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1715_ _1749_/D _1724_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
X_1577_ _1577_/B _1857_/A _1577_/A _1577_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XPHY_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput119 VPWR VGND pmatrix_row_out_n[2] _2090_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1500_ _1501_/S _1500_/A _1500_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
Xoutput108 VPWR VGND pmatrix_col_out_n[6] _1338_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput90 VPWR VGND pmatrix_col_out_n[19] _1384_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1362_ _1362_/X _1353_/D _1332_/X _1386_/B _1353_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1293_ _1435_/A _1311_/B _1311_/A _1423_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
X_1431_ _1431_/X _1430_/X _1367_/B _1429_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_23_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1629_ _1864_/A _1629_/X _1893_/A _1625_/X _1621_/A _1628_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a32o_2
XFILLER_36_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1980_ _1980_/Q fanout170/X _1980_/D _2042_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_0931_ _0934_/A _0949_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1414_ _1414_/X _1451_/A _1412_/Y _1471_/B _1413_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_2
X_1276_ VPWR VGND _1464_/A _1390_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1345_ VPWR VGND _1367_/B _1345_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout165 VPWR VGND fanout165/X fanout172/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout176 VPWR VGND fanout176/X fanout177/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout187 VPWR VGND _2066_/CLK _2065_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_10_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1130_ _1245_/B _1123_/X _1187_/B _1129_/X _1165_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_4
X_1061_ _1148_/D _0968_/X _0965_/X _1145_/A _1223_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1894_ _1621_/A _1893_/X _1892_/X _1894_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1963_ VGND VPWR _1963_/S input5/X _2067_/Q _1964_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_0914_ _0957_/B _1003_/B _2067_/Q _0914_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1259_ _1259_/B _1259_/X _1259_/A _1259_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1328_ _1423_/A _1328_/Y _1749_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_2093_ VGND VPWR _2093_/X _2093_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1113_ _1970_/Q _1154_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1044_ VPWR VGND _1044_/X _1036_/Y _1103_/B _1103_/A _1044_/B VGND VPWR sky130_fd_sc_hd__and4b_2
X_1877_ _1923_/B _1877_/Y _1877_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1946_ VGND VPWR _2059_/D _1946_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_28_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1800_ VGND VPWR _1996_/D _1800_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1662_ _2023_/Q _1664_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1731_ _1732_/A _1747_/B _1731_/A _1733_/A _1749_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
X_1593_ _1597_/S _1592_/X _2014_/Q _1552_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_2076_ VGND VPWR _2076_/X _2076_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1027_ _1103_/A _1025_/X _1148_/B _1023_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
XFILLER_38_155 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1929_ VGND VPWR _1929_/S _2023_/D _2021_/D _1929_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1645_ _1915_/A _1645_/Y _2019_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1576_ _1839_/A _1836_/A _1577_/C _2011_/Q _1836_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1714_ _1749_/D _1269_/B _1267_/X _1266_/X _1975_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__o31a_4
XPHY_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2059_ _2059_/Q fanout167/X _2059_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_59 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_103 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1430_ _1430_/X _1423_/A _1366_/X _1731_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
Xoutput109 VPWR VGND pmatrix_col_out_n[7] _1342_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput80 VPWR VGND pmatrix_col_out_n[0] _1296_/Y VGND VPWR sky130_fd_sc_hd__buf_4
X_1361_ _1361_/X _1386_/B _1324_/X _1353_/D _1353_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
Xoutput91 VPWR VGND pmatrix_col_out_n[1] _1310_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1292_ _1311_/B _1109_/B _1287_/Y _1290_/X _1288_/Y _1291_/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__o2111a_4
X_1559_ _1864_/A _1559_/Y _1526_/X _1893_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1628_ _2064_/Q _1628_/X _1626_/Y _1619_/B _1869_/B _1627_/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__a32o_2
XFILLER_36_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_301 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_143 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_165 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0930_ _1793_/S _0934_/A _1003_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_47_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1413_ _1413_/Y _1469_/A _1446_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_3_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1275_ VPWR VGND _2096_/A _1747_/B VGND VPWR sky130_fd_sc_hd__buf_2
X_1344_ _1344_/B _1345_/A _1350_/B _1344_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
Xfanout166 VPWR VGND fanout166/X fanout172/X VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout177 VPWR VGND fanout177/X fanout178/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout188 VPWR VGND _2065_/CLK _2063_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_8_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1060_ _1055_/Y _1058_/X _1221_/B _1059_/X _1066_/C _1056_/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__a221o_4
XFILLER_18_253 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1962_ VGND VPWR _2066_/D _1962_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_289 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1893_ _1893_/A _1893_/X _1893_/B _1621_/A _1897_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4bb_2
X_0913_ _2066_/Q _0914_/C _2065_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1327_ VPWR VGND _1423_/A _1394_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_1258_ _1259_/A _1259_/C _1259_/B _1258_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1189_ _1203_/A _1203_/B _1190_/C _1193_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_30_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2092_ VGND VPWR _2092_/X _2092_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1043_ VGND VPWR _1992_/Q _1956_/B _1991_/Q _1103_/B _1156_/B VGND VPWR sky130_fd_sc_hd__and4bb_2
X_1112_ VGND VPWR _1969_/D _1112_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_94 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1945_ VGND VPWR _1956_/D _1971_/D _2059_/Q _1946_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1876_ _2033_/Q _1831_/B _2033_/D _1875_/X _1874_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1730_ VGND VPWR _2088_/A _1730_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1661_ _1664_/C _2022_/Q _2020_/Q _2021_/Q _1671_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__and4_2
XFILLER_11_270 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1592_ _2014_/Q _2061_/Q _1552_/S _1592_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_2075_ VGND VPWR _2075_/X _2075_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1026_ _1233_/C _1103_/A _1157_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1928_ _1928_/B _1928_/X _2019_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1859_ _1859_/X _1915_/C _2009_/D _1870_/D VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_55_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1713_ VPWR VGND _2076_/A _1713_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1644_ _1915_/A _1870_/A _1644_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1575_ _1612_/B _1836_/B _1577_/B _1836_/C _1839_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
XPHY_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2058_ _2058_/Q fanout168/X _2058_/D _2060_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_1009_ _1963_/S _1956_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_32_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput70 VPWR VGND nmatrix_rowon_out_n[3] _2077_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_70 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1360_ VGND VPWR _1360_/X _1360_/A VGND VPWR sky130_fd_sc_hd__buf_1
Xoutput92 VPWR VGND pmatrix_col_out_n[20] _1385_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput81 VPWR VGND pmatrix_col_out_n[10] _1360_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1291_ _1290_/A _1290_/B _1290_/C _1291_/Y _1281_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__o211ai_2
X_1489_ _1489_/X _2006_/Q _1904_/A _2053_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1558_ _2054_/Q _1558_/Y _1557_/Y _1556_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1627_ _1621_/A _1627_/Y _1869_/B _2017_/Q _1893_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_2
XFILLER_39_273 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1412_ _1412_/Y _1435_/B _1412_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1343_ _1343_/Y _1343_/A _1457_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_51_213 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1274_ _1976_/D _1273_/X _1747_/B _2104_/A _1216_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
XFILLER_22_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_0989_ _0989_/B _0990_/D _1262_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
Xfanout167 VPWR VGND fanout167/X fanout172/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout189 VPWR VGND _2067_/CLK _2063_/CLK VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout178 VPWR VGND fanout178/X input9/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_221 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1892_ VGND VPWR _1897_/A _1610_/Y _1893_/A _1892_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1961_ VGND VPWR _1963_/S input4/X _2066_/Q _1962_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_0912_ _0957_/B _2046_/Q _0955_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1326_ _1412_/B _1394_/B _1435_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_24_246 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1257_ _1975_/Q _1259_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1188_ _1203_/B _1188_/B _1227_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_47_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_2091_ VGND VPWR _2091_/X _2091_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1042_ _1177_/B _1156_/B _1123_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1111_ VPWR VGND _1956_/B _1112_/A _1111_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_1875_ _1906_/A _1906_/C _2008_/D _1875_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1944_ VGND VPWR _2058_/D _1944_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1309_ _1309_/Y _1408_/A _1343_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_12_216 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_227 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1660_ _1660_/B _2022_/D _1784_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1591_ _1605_/A _2062_/Q _2015_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1025_ _1233_/A _1150_/B _1025_/X _1150_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_2074_ VGND VPWR _2074_/X _2074_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1927_ _2041_/D _1926_/X _1925_/X _1923_/X _1924_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1858_ _1858_/A _1915_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1789_ VGND VPWR _1793_/S _1992_/Q _1991_/Q _1790_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_113 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1643_ _1893_/B _1643_/Y _1665_/A _1913_/B _1913_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o31ai_2
X_1712_ _1744_/B _1713_/A _2081_/A _1712_/C VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
XANTENNA_1 _1411_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1574_ _1839_/A _1571_/X _1577_/A _1524_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21bo_2
XPHY_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2057_ _2057_/Q fanout167/X _2057_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _2105_/A _1963_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
Xoutput71 VPWR VGND nmatrix_rowon_out_n[4] _2078_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput93 VPWR VGND pmatrix_col_out_n[21] _1388_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput82 VPWR VGND pmatrix_col_out_n[11] _1361_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput60 VPWR VGND nmatrix_row_out_n[8] _1271_/X VGND VPWR sky130_fd_sc_hd__buf_4
X_1290_ _1290_/C _1290_/A _1290_/X _1290_/B _1290_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1626_ _1626_/A _1626_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_2
X_1557_ _1557_/B _1557_/Y _2007_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1488_ VPWR VGND _1904_/A _1665_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_22_163 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1342_ _1342_/X _1328_/Y _1460_/B _1341_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1411_ _1469_/A _1471_/B _1408_/Y _1411_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1273_ VGND VPWR _2104_/A _1273_/X _1216_/S _1976_/Q VGND VPWR sky130_fd_sc_hd__and3b_2
X_0988_ _1145_/B _1144_/A _0989_/B _0988_/B _1150_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1609_ VPWR VGND _1621_/A _2063_/Q VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout179 VPWR VGND _2034_/CLK fanout186/X VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout168 VPWR VGND fanout168/X fanout172/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_47_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1891_ _2036_/D _1890_/X _1889_/X _1887_/X _1888_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_0911_ _2044_/Q _0955_/B _2045_/Q _2043_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1960_ VGND VPWR _2065_/D _1960_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_52_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1325_ VPWR VGND _1435_/B _1355_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1256_ VGND VPWR _1267_/B _1252_/X _1253_/X _1259_/C _1255_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_2
X_1187_ _1203_/A _1245_/B _1187_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_47_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1110_ VGND VPWR _1110_/S _1109_/X _1969_/Q _1111_/B VGND VPWR sky130_fd_sc_hd__mux2_1
X_2090_ VGND VPWR _2090_/X _2090_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_21_206 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1041_ _1967_/Q _1041_/B _1148_/A _1066_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or3b_4
X_1874_ _1874_/X _1849_/X _2016_/D _1873_/X _1861_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
X_1943_ VGND VPWR _1977_/D _1970_/D _1836_/C _1944_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1308_ VPWR VGND _1343_/A _1446_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_1239_ _1290_/A _1220_/A _1093_/X _1029_/X _1166_/A _1138_/A VPWR VGND VGND VPWR
+ sky130_fd_sc_hd__o2111a_4
XFILLER_55_180 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
X_1590_ _1621_/D _2062_/Q _2015_/Q _1590_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__or3b_2
XFILLER_50_70 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_309 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1024_ VGND VPWR _1150_/C _1123_/A _1144_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
X_1926_ _2041_/Q _1819_/A _1926_/X _2016_/D _1882_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1857_ _1915_/B _1857_/Y _1857_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1788_ _1990_/D _1977_/D _1963_/S _0949_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_30_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_279 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1642_ _1913_/B _1641_/X _2018_/Q _1624_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1711_ _1712_/C _1376_/A _1717_/B _1717_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
XANTENNA_2 _1333_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_1573_ _1572_/Y _1867_/A _1513_/S _1839_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2056_ _2056_/Q fanout177/X _2056_/D _2063_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1007_ _1007_/Y _1007_/A _1259_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1909_ _2018_/D _1878_/B _1909_/X _2020_/D _1906_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_41_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput61 VPWR VGND nmatrix_row_out_n[9] _2082_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput72 VPWR VGND nmatrix_rowon_out_n[5] _2079_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput83 VPWR VGND pmatrix_col_out_n[12] _1362_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput50 VPWR VGND nmatrix_row_out_n[13] _2086_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput94 VPWR VGND pmatrix_col_out_n[22] _1392_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1556_ _2007_/Q _1556_/X _1870_/A _1557_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__and3_2
X_1625_ _1625_/X _1624_/X _1633_/B _1870_/A _1869_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a31o_2
X_1487_ VPWR VGND _1665_/A _1870_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_39_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_2039_ _2039_/Q fanout166/X _2039_/D _2039_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_9_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1410_ _1409_/Y _1408_/Y _1400_/X _1471_/B _1410_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__o211a_2
X_1272_ VPWR VGND _1747_/B _1749_/C VGND VPWR sky130_fd_sc_hd__buf_6
X_1341_ _1341_/Y _1408_/B _1457_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_0987_ _1150_/B _1177_/B _1126_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__or2_4
X_1608_ _1897_/A _1608_/X _1607_/Y _1893_/A _1836_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__o22a_2
X_1539_ _1539_/B _1539_/Y _1893_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
Xfanout169 VPWR VGND fanout169/X fanout171/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_47_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_270 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_234 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1890_ _2036_/Q _1831_/B _1890_/X _1836_/C _1882_/Y VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_0910_ _1993_/Q _1994_/Q _1003_/A _1992_/Q _1991_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4_2
XFILLER_45_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1324_ VPWR VGND _1324_/X _1324_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1255_ VGND VPWR _1255_/X _1081_/Y _1198_/Y _1066_/A _1066_/C _1066_/D VGND VPWR
+ sky130_fd_sc_hd__a311o_2
X_1186_ _1190_/A _1190_/B _1193_/B _1193_/A _1185_/X _1318_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111ai_4
X_1040_ _1044_/B _1036_/Y _1040_/D _1041_/B _1037_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__and4bb_4
X_1942_ VGND VPWR _2057_/D _1942_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1873_ _1873_/X _1906_/D _2012_/D _2014_/D _1878_/B VGND VPWR _1872_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_28_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_329 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1307_ _1307_/Y _1451_/A _1471_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__nand2_2
X_1169_ _1169_/A _1350_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_8
X_1238_ _1262_/B _1262_/C _1238_/X _1238_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_18_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1023_ _1023_/B _1023_/X _1262_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
X_1925_ _2018_/D _1915_/B _1925_/X _1928_/B _1858_/A _2020_/D VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
X_1787_ VGND VPWR _1989_/D _1787_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_1856_ _1889_/B _1856_/Y _1877_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_29_104 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_107 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_203 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_85 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_321 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1572_ _2057_/Q _1572_/Y _2010_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1641_ _1621_/A _1893_/A _2017_/Q _2064_/Q _2018_/Q _1641_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111a_2
X_1710_ VPWR VGND _2075_/A _1710_/A VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA_3 _1414_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_2055_ _2055_/Q fanout173/X _2055_/D _2066_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1006_ VPWR VGND _1216_/S _1259_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_1908_ _2038_/D _1907_/X _1903_/Y _1905_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a21o_2
X_1839_ _1839_/A _1923_/B _1839_/X _1839_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_9_317 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput73 VPWR VGND nmatrix_rowon_out_n[6] _2080_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput95 VPWR VGND pmatrix_col_out_n[23] _1393_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput40 VPWR VGND nmatrix_col_out_n[3] _1421_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput84 VPWR VGND pmatrix_col_out_n[13] _1365_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput51 VPWR VGND nmatrix_row_out_n[14] _2087_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput62 VPWR VGND nmatrix_rowon_out_n[0] _2074_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1624_ VPWR VGND _2064_/Q _1624_/X _2017_/Q VGND VPWR sky130_fd_sc_hd__and2_2
X_1555_ VPWR VGND _2014_/D _1555_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_1486_ VPWR VGND _1870_/A _1977_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_2038_ _2038_/Q fanout166/X _2038_/D _2039_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_6_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_125 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_169 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_72 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1340_ _1457_/C _1435_/A _1471_/A VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_4
X_1271_ VPWR VGND _1271_/X _1729_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_235 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_0986_ VPWR VGND _1126_/A _2001_/Q VGND VPWR sky130_fd_sc_hd__buf_6
X_1607_ _1612_/B _1897_/A _1893_/A _1607_/Y VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1538_ _2059_/Q _1538_/B _1539_/B _1538_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
X_1469_ _1469_/A _1749_/A _1469_/X _1469_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__or3_2
XFILLER_47_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_282 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1323_ _1404_/C _1324_/A _1435_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_38_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1185_ _1198_/A _1226_/B _1289_/A _1185_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1254_ _1212_/B _1173_/B _1252_/X _1267_/B _1212_/A VPWR VGND VGND VPWR sky130_fd_sc_hd__a211oi_2
X_0969_ _1991_/Q _1993_/Q _1992_/Q _2105_/A _1122_/B VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_30_208 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_65 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
X_1872_ _1872_/X _1865_/X _1870_/D _1868_/Y _1871_/X VGND VPWR VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_21_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1941_ VGND VPWR _1977_/D _1969_/D _1870_/C _1942_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_1306_ VPWR VGND _1451_/A _1399_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_1237_ _1222_/X _1264_/A _1235_/Y _1242_/B VGND VPWR VGND VPWR sky130_fd_sc_hd__a21oi_2
X_1168_ VPWR VGND _1317_/A _1169_/A _1317_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_44_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
X_1099_ _1238_/C _1098_/X _1019_/X _1020_/X _1104_/A _1099_/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o32a_2
XFILLER_20_263 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_1022_ _2105_/A _1991_/Q _1023_/B _1993_/Q _1992_/Q VPWR VGND VGND VPWR sky130_fd_sc_hd__or4b_2
X_1855_ _2031_/Q _1831_/B _2031_/D _1854_/X _1853_/X VPWR VGND VGND VPWR sky130_fd_sc_hd__a22o_2
X_1924_ _1849_/X _1924_/Y _1670_/B _1784_/S VGND VPWR VGND VPWR sky130_fd_sc_hd__o21ai_2
X_1786_ VGND VPWR _1786_/S _1989_/Q input8/X _1787_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1571_ _1836_/C _1596_/A _1571_/X _2011_/Q _1621_/D VPWR VGND VGND VPWR sky130_fd_sc_hd__or4_2
X_1640_ _1632_/B _1606_/A _2017_/Q _2064_/Q _2018_/Q _1913_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o2111a_2
XANTENNA_4 _1415_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_2054_ _2054_/Q fanout167/X _2054_/D _2059_/CLK VGND VPWR VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_1005_ VPWR VGND _1259_/B _1110_/S VGND VPWR sky130_fd_sc_hd__buf_6
X_1907_ _1907_/X _1882_/Y _2038_/Q _2013_/D _1819_/A VGND VPWR _1906_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_1838_ _1524_/B _1524_/A _1915_/A _1839_/C VGND VPWR VGND VPWR sky130_fd_sc_hd__o21a_2
X_1769_ VPWR VGND _1982_/Q _1775_/C _1769_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_25_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput52 VPWR VGND nmatrix_row_out_n[15] _2088_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput41 VPWR VGND nmatrix_col_out_n[4] _1422_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput30 VPWR VGND nmatrix_col_out_n[23] _1459_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput63 VPWR VGND nmatrix_rowon_out_n[10] _2084_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput74 VPWR VGND nmatrix_rowon_out_n[7] _2081_/X VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput85 VPWR VGND pmatrix_col_out_n[14] _1369_/Y VGND VPWR sky130_fd_sc_hd__buf_4
Xoutput96 VPWR VGND pmatrix_col_out_n[24] _1395_/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_48_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_1485_ VGND VPWR _1869_/B _1557_/B _2053_/Q _1485_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_1623_ _2017_/Q _1633_/B _2064_/Q VGND VPWR VGND VPWR sky130_fd_sc_hd__nor2_2
X_1554_ _2061_/Q _2014_/Q _1555_/A _1550_/X _1553_/X _1864_/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hd__o221a_2
.ends

